CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
7 74LS251
144 923 1135 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
5130 0 0
2
45434.7 0
0
7 74LS251
144 1082 1066 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
391 0 0
2
45434.7 0
0
7 74LS251
144 928 914 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
3124 0 0
2
45434.7 0
0
7 74LS251
144 1003 796 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
3421 0 0
2
45434.7 0
0
7 74LS251
144 590 503 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U7
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
8157 0 0
2
45434.7 0
0
7 74LS251
144 592 397 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
5572 0 0
2
45434.7 0
0
7 74LS251
144 591 294 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
8901 0 0
2
45434.7 0
0
7 74LS251
144 592 191 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
7361 0 0
2
45434.7 0
0
8 Hex Key~
166 1112 35 0 11 12
0 11 13 15 16 0 0 0 0 0
8 56
0
0 0 4640 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4747 0 0
2
45434.6 0
0
7 74LS251
144 588 96 0 1 29
0 0
0
0 0 4832 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 0 0 0 0 0
1 U
972 0 0
2
45434.6 0
0
12 Hex Display~
7 492 48 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3472 0 0
2
45434.6 0
0
6 74136~
219 460 824 0 3 22
0 3 6 2
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9998 0 0
2
45434.6 0
0
6 74136~
219 406 751 0 3 22
0 4 7 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3536 0 0
2
45434.6 0
0
6 74136~
219 351 661 0 3 22
0 5 8 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4597 0 0
2
45434.6 0
0
6 74136~
219 300 579 0 3 22
0 10 9 5
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3835 0 0
2
45434.6 0
0
6 74136~
219 246 457 0 3 22
0 12 11 10
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3670 0 0
2
45434.6 0
0
6 74136~
219 195 371 0 3 22
0 14 13 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5616 0 0
2
45434.6 0
0
8 Hex Key~
166 58 50 0 11 12
0 11 13 15 16 0 0 0 0 0
8 56
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9323 0 0
2
45434.6 0
0
6 74136~
219 90 203 0 3 22
0 15 16 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
317 0 0
2
45434.6 0
0
12 Hex Display~
7 410 62 0 18 19
10 10 12 14 16 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3108 0 0
2
45434.6 0
0
6 74136~
219 141 266 0 3 22
0 17 15 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4299 0 0
2
45434.6 0
0
8 Hex Key~
166 238 536 0 11 12
0 6 7 8 9 0 0 0 0 0
8 56
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9672 0 0
2
45434.6 0
0
33
1 11 0 0 0 0 0 9 7 0 0 3
1121 59
1121 285
623 285
10 2 0 0 0 0 0 7 9 0 0 3
623 276
1115 276
1115 59
3 9 0 0 0 0 0 9 7 0 0 3
1109 59
1109 267
623 267
11 1 0 0 0 0 0 8 9 0 0 3
624 182
1121 182
1121 59
2 10 0 0 0 0 0 9 8 0 0 3
1115 59
1115 173
624 173
9 3 0 0 0 0 0 8 9 0 0 3
624 164
1109 164
1109 59
3 9 0 0 0 0 0 9 10 0 0 3
1109 59
1109 69
620 69
2 10 0 0 0 0 0 9 10 0 0 3
1115 59
1115 78
620 78
1 11 0 0 0 0 0 9 10 0 0 3
1121 59
1121 87
620 87
3 1 2 0 0 8320 0 12 11 0 0 3
493 824
501 824
501 72
3 2 3 0 0 8320 0 13 11 0 0 3
439 751
495 751
495 72
3 3 4 0 0 8320 0 14 11 0 0 3
384 661
489 661
489 72
3 4 5 0 0 4224 0 15 11 0 0 3
333 579
483 579
483 72
2 1 6 0 0 8320 0 12 22 0 0 3
444 833
247 833
247 560
3 1 3 0 0 0 0 13 12 0 0 3
439 751
439 815
444 815
2 2 7 0 0 4224 0 22 13 0 0 3
241 560
241 760
390 760
2 3 8 0 0 8320 0 14 22 0 0 3
335 670
235 670
235 560
3 1 4 0 0 0 0 14 13 0 0 4
384 661
388 661
388 742
390 742
3 1 5 0 0 0 0 15 14 0 0 4
333 579
332 579
332 652
335 652
4 2 9 0 0 8320 0 22 15 0 0 3
229 560
229 588
284 588
3 1 10 0 0 8192 0 16 15 0 0 4
279 457
281 457
281 570
284 570
3 1 10 0 0 4224 0 16 20 0 0 3
279 457
419 457
419 86
2 1 11 0 0 8320 0 16 18 0 0 3
230 466
67 466
67 74
3 1 12 0 0 8192 0 17 16 0 0 4
228 371
229 371
229 448
230 448
3 2 12 0 0 4224 0 17 20 0 0 3
228 371
413 371
413 86
2 2 13 0 0 4224 0 18 17 0 0 3
61 74
61 380
179 380
3 1 14 0 0 8192 0 21 17 0 0 4
174 266
176 266
176 362
179 362
3 3 14 0 0 4224 0 21 20 0 0 3
174 266
407 266
407 86
3 2 15 0 0 4224 0 18 21 0 0 3
55 74
55 275
125 275
3 1 15 0 0 0 0 18 19 0 0 3
55 74
55 194
74 194
4 2 16 0 0 4096 0 18 19 0 0 3
49 74
49 212
74 212
4 4 16 0 0 8320 0 18 20 0 0 4
49 74
49 173
401 173
401 86
3 1 17 0 0 8320 0 19 21 0 0 4
123 203
122 203
122 257
125 257
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
