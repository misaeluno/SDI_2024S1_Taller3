CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 2070 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
96
8 Hex Key~
166 17 3333 0 11 12
0 31 23 24 21 0 0 0 0 0
2 50
0
0 0 4640 180
0
4 KPD5
20 -2 48 6
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5130 0 0
2
45438.8 0
0
13 Logic Switch~
5 1726 155 0 1 11
0 15
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
45438.8 0
0
13 Logic Switch~
5 1160 22 0 1 11
0 91
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
45438.8 1
0
7 Buffer~
58 865 1220 0 2 22
0 6 3
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35C
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 30 0
1 U
3421 0 0
2
45438.8 0
0
7 Buffer~
58 802 1221 0 2 22
0 7 4
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35B
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 30 0
1 U
8157 0 0
2
45438.8 0
0
7 Buffer~
58 746 1213 0 2 22
0 8 5
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35A
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 30 0
1 U
5572 0 0
2
45438.8 0
0
7 Ground~
168 1653 13 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
45438.8 0
0
9 CC 7-Seg~
183 1653 91 0 16 19
10 18 17 16 14 13 12 11 15 2
1 1 1 1 0 1 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
7361 0 0
2
45438.8 0
0
9 Inverter~
13 129 1840 0 2 22
0 21 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U29A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 24 0
1 U
4747 0 0
2
45438.8 0
0
9 Inverter~
13 210 1741 0 2 22
0 23 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U27A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
972 0 0
2
45438.8 0
0
9 Inverter~
13 157 1750 0 2 22
0 24 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U21A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
3472 0 0
2
45438.8 0
0
9 Inverter~
13 110 1759 0 2 22
0 21 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 29 0
1 U
9998 0 0
2
45438.8 0
0
9 2-In AND~
219 215 1831 0 3 22
0 24 22 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
3536 0 0
2
45438.8 0
0
5 7415~
219 273 1750 0 4 22
0 25 26 27 28
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 12 0
1 U
4597 0 0
2
45438.8 0
0
8 2-In OR~
219 533 1759 0 3 22
0 28 29 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
3835 0 0
2
45438.8 0
0
9 Inverter~
13 203 1325 0 2 22
0 24 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 29 0
1 U
3670 0 0
2
45438.8 0
0
9 2-In AND~
219 326 947 0 3 22
0 21 23 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
5616 0 0
2
45438.8 0
0
9 Inverter~
13 120 1009 0 2 22
0 21 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 29 0
1 U
9323 0 0
2
5.90125e-315 0
0
9 Inverter~
13 163 1000 0 2 22
0 24 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 29 0
1 U
317 0 0
2
5.90125e-315 0
0
9 Inverter~
13 203 991 0 2 22
0 23 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 29 0
1 U
3108 0 0
2
5.90125e-315 0
0
5 7415~
219 349 1000 0 4 22
0 36 35 34 33
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 8 0
1 U
4299 0 0
2
5.90125e-315 0
0
9 Inverter~
13 215 2268 0 2 22
0 24 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 27 0
1 U
9672 0 0
2
5.90125e-315 0
0
9 Inverter~
13 206 2215 0 2 22
0 23 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 27 0
1 U
7876 0 0
2
5.90125e-315 0
0
9 Inverter~
13 220 2172 0 2 22
0 21 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 27 0
1 U
6369 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 402 2259 0 3 22
0 23 37 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
9172 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 345 2224 0 3 22
0 38 24 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
7100 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 394 2181 0 3 22
0 39 24 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
3820 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 562 2173 0 5 22
0 31 42 41 40 6
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 25 0
1 U
7678 0 0
2
5.90125e-315 0
0
9 Inverter~
13 233 2079 0 2 22
0 24 45
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 27 0
1 U
961 0 0
2
5.90125e-315 0
0
9 Inverter~
13 233 2027 0 2 22
0 21 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 27 0
1 U
3178 0 0
2
5.90125e-315 0
0
9 Inverter~
13 201 1973 0 2 22
0 24 49
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 27 0
1 U
3409 0 0
2
5.90125e-315 0
0
9 Inverter~
13 144 1991 0 2 22
0 21 48
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28F
-14 -18 14 -10
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 23 0
1 U
3951 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 371 2070 0 3 22
0 23 45 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
8885 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 367 2018 0 3 22
0 23 46 44
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
3780 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 309 1982 0 3 22
0 49 48 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
9265 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 554 1976 0 5 22
0 31 47 44 43 7
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 25 0
1 U
9442 0 0
2
5.90125e-315 0
0
9 Inverter~
13 142 1685 0 2 22
0 21 50
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 21 0
1 U
9424 0 0
2
5.90125e-315 0
0
9 Inverter~
13 198 1667 0 2 22
0 31 51
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 20 0
1 U
9968 0 0
2
5.90125e-315 0
0
9 Inverter~
13 167 1622 0 2 22
0 23 52
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 20 0
1 U
9281 0 0
2
5.90125e-315 0
0
9 Inverter~
13 90 1613 0 2 22
0 31 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 20 0
1 U
8464 0 0
2
5.90125e-315 0
0
9 Inverter~
13 250 1577 0 2 22
0 24 57
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 20 0
1 U
7168 0 0
2
5.90125e-315 0
0
9 Inverter~
13 171 1568 0 2 22
0 23 58
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 20 0
1 U
3171 0 0
2
5.90125e-315 0
0
9 Inverter~
13 221 1534 0 2 22
0 24 60
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 20 0
1 U
4139 0 0
2
5.90125e-315 0
0
8 Hex Key~
166 55 2304 0 11 12
0 31 23 24 21 0 0 0 0 0
2 50
0
0 0 4656 180
0
4 KPD4
20 -2 48 6
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6435 0 0
2
5.90125e-315 0
0
9 Inverter~
13 182 1506 0 2 22
0 21 62
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 14 0
1 U
5283 0 0
2
5.90125e-315 0
0
9 Inverter~
13 231 1497 0 2 22
0 24 63
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 14 0
1 U
6874 0 0
2
5.90125e-315 0
0
9 Inverter~
13 278 1488 0 2 22
0 23 64
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 14 0
1 U
5305 0 0
2
5.90125e-315 0
0
5 7415~
219 365 1676 0 4 22
0 51 24 50 54
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 19 0
1 U
34 0 0
2
5.90125e-315 0
0
5 7415~
219 366 1568 0 4 22
0 31 58 57 56
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 19 0
1 U
969 0 0
2
5.90125e-315 0
0
5 7415~
219 323 1534 0 4 22
0 23 60 21 59
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 19 0
1 U
8402 0 0
2
5.90125e-315 0
0
5 7415~
219 323 1622 0 4 22
0 53 52 24 55
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 15 0
1 U
3751 0 0
2
5.90125e-315 0
0
5 7415~
219 363 1497 0 4 22
0 64 63 62 61
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 15 0
1 U
4292 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 524 1528 0 3 22
0 66 65 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
6118 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 433 1646 0 3 22
0 55 54 65
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
34 0 0
2
5.90125e-315 0
0
8 3-In OR~
219 423 1506 0 4 22
0 61 59 56 66
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U22A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 17 0
1 U
6357 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 533 1320 0 5 22
0 31 23 30 21 10
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
319 0 0
2
5.90125e-315 0
0
9 Inverter~
13 198 1229 0 2 22
0 24 68
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
3976 0 0
2
5.90125e-315 0
0
9 Inverter~
13 160 1211 0 2 22
0 21 69
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
7634 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 384 1220 0 3 22
0 69 68 67
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
523 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 311 1194 0 3 22
0 24 21 70
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
6748 0 0
2
5.90125e-315 0
0
9 Inverter~
13 97 1170 0 2 22
0 23 71
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
6901 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 568 1174 0 5 22
0 31 71 70 67 19
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
842 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 575 1078 0 5 22
0 32 33 24 31 20
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
3277 0 0
2
45438.8 3
0
6 74136~
219 127 769 0 3 22
0 24 21 73
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4212 0 0
2
45438.8 5
0
6 74136~
219 129 719 0 3 22
0 23 24 74
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
4720 0 0
2
45438.8 6
0
6 74136~
219 127 667 0 3 22
0 31 23 75
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5551 0 0
2
45438.8 7
0
6 74136~
219 126 612 0 3 22
0 80 31 79
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6986 0 0
2
45438.8 8
0
6 74136~
219 133 564 0 3 22
0 84 80 81
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
8745 0 0
2
45438.8 9
0
6 74136~
219 126 513 0 3 22
0 85 84 82
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9592 0 0
2
45438.8 10
0
6 74136~
219 200 448 0 3 22
0 72 85 83
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8748 0 0
2
45438.8 11
0
14 Logic Display~
6 1417 34 0 1 2
10 90
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90125e-315 0
0
14 Logic Display~
6 1382 24 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.90125e-315 5.26354e-315
0
14 Logic Display~
6 1354 23 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
5.90125e-315 5.30499e-315
0
14 Logic Display~
6 1332 23 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
5.90125e-315 5.32571e-315
0
14 Logic Display~
6 1298 27 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
5.90125e-315 5.34643e-315
0
14 Logic Display~
6 1273 31 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.90125e-315 5.3568e-315
0
14 Logic Display~
6 1250 33 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.90125e-315 5.36716e-315
0
14 Logic Display~
6 1215 34 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6263 0 0
2
5.90125e-315 5.37752e-315
0
6 74136~
219 385 355 0 3 22
0 77 21 76
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4900 0 0
2
5.90125e-315 5.38788e-315
0
6 74136~
219 335 331 0 3 22
0 78 24 77
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8783 0 0
2
5.90125e-315 5.39306e-315
0
6 74136~
219 284 295 0 3 22
0 86 23 78
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3221 0 0
2
5.90125e-315 5.39824e-315
0
6 74136~
219 237 266 0 3 22
0 87 31 86
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3215 0 0
2
5.90125e-315 5.40342e-315
0
6 74136~
219 186 225 0 3 22
0 88 80 87
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7903 0 0
2
5.90125e-315 5.4086e-315
0
7 74LS251
144 1023 801 0 14 29
0 96 97 98 99 100 76 101 73 92
93 94 91 102 90
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7121 0 0
2
45438.8 12
0
7 74LS251
144 1027 699 0 14 29
0 103 104 105 106 107 77 3 74 92
93 94 91 108 11
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4484 0 0
2
45438.8 13
0
7 74LS251
144 1027 599 0 14 29
0 109 110 111 112 113 78 4 75 92
93 94 91 114 12
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5996 0 0
2
45438.8 14
0
7 74LS251
144 1027 492 0 14 29
0 115 116 117 118 119 86 5 79 92
93 94 91 120 13
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7804 0 0
2
45438.8 15
0
7 74LS251
144 1028 389 0 14 29
0 121 122 123 124 125 87 9 81 92
93 94 91 126 14
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5523 0 0
2
45438.8 16
0
7 74LS251
144 1034 287 0 14 29
0 127 128 129 130 131 88 10 82 92
93 94 91 132 16
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3330 0 0
2
45438.8 17
0
7 74LS251
144 1033 187 0 14 29
0 133 134 135 136 137 89 19 83 92
93 94 91 138 17
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3465 0 0
2
45438.8 18
0
8 Hex Key~
166 1115 33 0 11 12
0 94 93 92 139 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8396 0 0
2
45438.8 19
0
7 74LS251
144 1033 94 0 14 29
0 140 141 142 143 144 72 20 72 92
93 94 91 145 18
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3685 0 0
2
45438.8 20
0
8 Hex Key~
166 15 40 0 11 12
0 80 84 85 72 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7849 0 0
2
45438.8 22
0
6 74136~
219 89 163 0 3 22
0 85 72 89
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6343 0 0
2
45438.8 23
0
6 74136~
219 138 193 0 3 22
0 89 84 88
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7376 0 0
2
45438.8 25
0
8 Hex Key~
166 52 42 0 11 12
0 21 24 23 31 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9156 0 0
2
45438.8 26
0
209
4 1 0 0 0 0 0 1 93 0 0 2
24 3309
24 64
2 3 0 0 0 0 0 93 1 0 0 2
18 64
18 3309
2 3 0 0 0 0 0 1 93 0 0 2
12 3309
12 64
4 1 0 0 0 0 0 93 1 0 0 2
6 64
6 3309
2 7 3 0 0 4224 0 4 85 0 0 3
865 1205
865 726
995 726
7 2 4 0 0 8320 0 86 5 0 0 3
995 626
802 626
802 1206
2 7 5 0 0 4224 0 6 87 0 0 3
746 1198
746 519
995 519
1 5 6 0 0 4224 0 4 28 0 0 3
865 1235
865 2173
595 2173
5 1 7 0 0 8320 0 36 5 0 0 3
587 1976
802 1976
802 1236
1 3 8 0 0 4224 0 6 15 0 0 3
746 1228
746 1759
566 1759
7 3 9 0 0 8320 0 88 53 0 0 6
996 416
710 416
710 1301
709 1301
709 1528
557 1528
7 5 10 0 0 8320 0 89 56 0 0 6
1002 314
696 314
696 1319
574 1319
574 1320
566 1320
14 7 11 0 0 8192 0 85 8 0 0 3
1059 735
1668 735
1668 127
6 14 12 0 0 8192 0 8 86 0 0 3
1662 127
1662 635
1059 635
14 5 13 0 0 4224 0 87 8 0 0 3
1059 528
1656 528
1656 127
4 14 14 0 0 8320 0 8 88 0 0 3
1650 127
1650 425
1060 425
1 8 15 0 0 4224 0 2 8 0 0 3
1712 155
1674 155
1674 127
14 3 16 0 0 4224 0 89 8 0 0 3
1066 323
1644 323
1644 127
2 14 17 0 0 8320 0 8 90 0 0 3
1638 127
1638 223
1065 223
14 1 18 0 0 4224 0 92 8 0 0 3
1065 130
1632 130
1632 127
5 7 19 0 0 8320 0 62 90 0 0 4
601 1174
682 1174
682 214
1001 214
5 7 20 0 0 8320 0 63 92 0 0 4
608 1078
664 1078
664 121
1001 121
9 1 2 0 0 4224 0 8 7 0 0 2
1653 49
1653 21
1 0 21 0 0 4096 0 9 0 0 102 2
114 1840
61 1840
2 2 22 0 0 4224 0 9 13 0 0 2
150 1840
191 1840
1 0 23 0 0 4096 0 10 0 0 104 2
195 1741
49 1741
1 0 24 0 0 4096 0 11 0 0 103 2
142 1750
55 1750
2 1 25 0 0 4224 0 10 14 0 0 2
231 1741
249 1741
2 2 26 0 0 4224 0 11 14 0 0 2
178 1750
249 1750
1 0 21 0 0 0 0 12 0 0 102 2
95 1759
61 1759
2 3 27 0 0 4224 0 12 14 0 0 2
131 1759
249 1759
4 1 28 0 0 4224 0 14 15 0 0 2
294 1750
520 1750
3 2 29 0 0 4224 0 13 15 0 0 4
236 1831
398 1831
398 1768
520 1768
1 0 24 0 0 4096 0 13 0 0 103 2
191 1822
55 1822
4 0 21 0 0 4096 0 56 0 0 102 2
516 1334
61 1334
1 0 24 0 0 0 0 16 0 0 103 2
188 1325
55 1325
2 3 30 0 0 4224 0 16 56 0 0 2
224 1325
516 1325
2 0 23 0 0 4096 0 56 0 0 104 2
516 1316
49 1316
1 0 31 0 0 4096 0 56 0 0 105 2
516 1307
43 1307
1 0 21 0 0 0 0 17 0 0 102 2
302 938
61 938
2 0 23 0 0 0 0 17 0 0 104 2
302 956
49 956
3 1 32 0 0 12416 0 17 63 0 0 4
347 947
433 947
433 1065
558 1065
4 0 31 0 0 4096 0 63 0 0 105 2
558 1092
43 1092
3 0 24 0 0 4096 0 63 0 0 103 2
558 1083
55 1083
2 4 33 0 0 4224 0 63 21 0 0 4
558 1074
378 1074
378 1000
370 1000
1 0 21 0 0 0 0 18 0 0 102 2
105 1009
61 1009
1 0 24 0 0 0 0 19 0 0 103 2
148 1000
55 1000
1 0 23 0 0 0 0 20 0 0 104 2
188 991
49 991
3 2 34 0 0 4224 0 21 18 0 0 2
325 1009
141 1009
2 2 35 0 0 4224 0 21 19 0 0 2
325 1000
184 1000
2 1 36 0 0 4224 0 20 21 0 0 2
224 991
325 991
1 0 23 0 0 0 0 25 0 0 104 2
378 2250
49 2250
1 0 24 0 0 0 0 22 0 0 103 2
200 2268
55 2268
2 2 37 0 0 4224 0 22 25 0 0 2
236 2268
378 2268
2 0 24 0 0 0 0 26 0 0 103 2
321 2233
55 2233
1 0 23 0 0 0 0 23 0 0 104 2
191 2215
49 2215
2 1 38 0 0 4224 0 23 26 0 0 2
227 2215
321 2215
2 0 24 0 0 0 0 27 0 0 103 2
370 2190
55 2190
1 0 21 0 0 0 0 24 0 0 102 2
205 2172
61 2172
2 1 39 0 0 4224 0 24 27 0 0 2
241 2172
370 2172
4 3 40 0 0 12416 0 28 25 0 0 4
545 2187
516 2187
516 2259
423 2259
3 3 41 0 0 12416 0 28 26 0 0 4
545 2178
470 2178
470 2224
366 2224
3 2 42 0 0 12416 0 27 28 0 0 4
415 2181
451 2181
451 2169
545 2169
1 0 31 0 0 0 0 28 0 0 105 2
545 2160
43 2160
3 4 43 0 0 4224 0 33 36 0 0 4
392 2070
529 2070
529 1990
537 1990
3 3 44 0 0 12416 0 34 36 0 0 4
388 2018
421 2018
421 1981
537 1981
1 0 24 0 0 0 0 29 0 0 103 2
218 2079
55 2079
1 0 23 0 0 0 0 34 0 0 104 2
343 2009
49 2009
2 2 45 0 0 4224 0 29 33 0 0 2
254 2079
347 2079
1 0 23 0 0 0 0 33 0 0 104 2
347 2061
49 2061
1 0 21 0 0 0 0 30 0 0 102 2
218 2027
61 2027
2 2 46 0 0 4224 0 30 34 0 0 2
254 2027
343 2027
3 2 47 0 0 12416 0 35 36 0 0 4
330 1982
381 1982
381 1972
537 1972
2 2 48 0 0 4224 0 35 32 0 0 2
285 1991
165 1991
2 1 49 0 0 4224 0 31 35 0 0 2
222 1973
285 1973
1 0 21 0 0 0 0 32 0 0 102 2
129 1991
61 1991
1 0 24 0 0 0 0 31 0 0 103 2
186 1973
55 1973
1 0 31 0 0 0 0 36 0 0 105 2
537 1963
43 1963
1 0 21 0 0 0 0 37 0 0 102 2
127 1685
61 1685
2 3 50 0 0 4224 0 37 48 0 0 2
163 1685
341 1685
2 0 24 0 0 0 0 48 0 0 103 2
341 1676
55 1676
1 0 31 0 0 0 0 38 0 0 105 2
183 1667
43 1667
2 1 51 0 0 4224 0 38 48 0 0 2
219 1667
341 1667
1 0 23 0 0 0 0 39 0 0 104 2
152 1622
49 1622
2 2 52 0 0 4224 0 39 51 0 0 2
188 1622
299 1622
1 0 31 0 0 0 0 40 0 0 105 2
75 1613
43 1613
2 1 53 0 0 4224 0 40 51 0 0 2
111 1613
299 1613
3 0 24 0 0 0 0 51 0 0 103 2
299 1631
55 1631
4 2 54 0 0 4224 0 48 54 0 0 4
386 1676
412 1676
412 1655
420 1655
4 1 55 0 0 4224 0 51 54 0 0 4
344 1622
412 1622
412 1637
420 1637
4 3 56 0 0 8320 0 49 55 0 0 4
387 1568
402 1568
402 1515
410 1515
1 0 24 0 0 0 0 41 0 0 103 2
235 1577
55 1577
1 0 23 0 0 0 0 42 0 0 104 2
156 1568
49 1568
2 3 57 0 0 4224 0 41 49 0 0 2
271 1577
342 1577
2 2 58 0 0 4224 0 42 49 0 0 2
192 1568
342 1568
1 0 31 0 0 0 0 49 0 0 105 2
342 1559
43 1559
3 0 21 0 0 0 0 50 0 0 102 2
299 1543
61 1543
1 0 24 0 0 0 0 43 0 0 103 2
206 1534
55 1534
4 2 59 0 0 4224 0 50 55 0 0 4
344 1534
381 1534
381 1506
411 1506
2 2 60 0 0 4224 0 43 50 0 0 2
242 1534
299 1534
0 1 23 0 0 0 0 0 50 104 0 2
49 1525
299 1525
1 4 21 0 0 4224 0 96 44 0 0 4
61 66
61 1840
62 1840
62 2280
2 3 24 0 0 4224 0 96 44 0 0 4
55 66
55 1822
56 1822
56 2280
3 2 23 0 0 4224 0 96 44 0 0 4
49 66
49 1741
50 1741
50 2280
4 1 31 0 0 4224 0 96 44 0 0 4
43 66
43 1307
44 1307
44 2280
4 1 61 0 0 4224 0 52 55 0 0 2
384 1497
410 1497
2 3 62 0 0 4224 0 45 52 0 0 2
203 1506
339 1506
2 2 63 0 0 4224 0 52 46 0 0 2
339 1497
252 1497
2 1 64 0 0 4224 0 47 52 0 0 2
299 1488
339 1488
1 1 21 0 0 0 0 96 45 0 0 3
61 66
61 1506
167 1506
2 1 24 0 0 0 0 96 46 0 0 3
55 66
55 1497
216 1497
3 1 23 0 0 0 0 96 47 0 0 3
49 66
49 1488
263 1488
2 3 65 0 0 8320 0 53 54 0 0 4
511 1537
490 1537
490 1646
466 1646
4 1 66 0 0 4224 0 55 53 0 0 4
456 1506
489 1506
489 1519
511 1519
3 4 67 0 0 12416 0 59 62 0 0 4
405 1220
471 1220
471 1188
551 1188
2 2 68 0 0 4224 0 59 57 0 0 2
360 1229
219 1229
2 1 69 0 0 4224 0 58 59 0 0 2
181 1211
360 1211
2 1 24 0 0 0 0 96 57 0 0 3
55 66
55 1229
183 1229
1 1 21 0 0 0 0 96 58 0 0 3
61 66
61 1211
145 1211
3 3 70 0 0 12416 0 60 62 0 0 4
332 1194
368 1194
368 1179
551 1179
1 2 21 0 0 0 0 96 60 0 0 3
61 66
61 1203
287 1203
2 1 24 0 0 0 0 96 60 0 0 3
55 66
55 1185
287 1185
2 2 71 0 0 4224 0 61 62 0 0 2
118 1170
551 1170
3 1 23 0 0 0 0 96 61 0 0 3
49 66
49 1170
82 1170
4 1 31 0 0 0 0 96 62 0 0 3
43 66
43 1161
551 1161
4 1 72 0 0 4096 0 93 70 0 0 3
6 64
6 439
184 439
3 8 73 0 0 4224 0 64 84 0 0 4
160 769
603 769
603 837
991 837
3 8 74 0 0 16512 0 65 85 0 0 5
162 719
162 724
577 724
577 735
995 735
3 8 75 0 0 12416 0 66 86 0 0 4
160 667
566 667
566 635
995 635
3 6 76 0 0 8320 0 79 84 0 0 4
418 355
528 355
528 819
991 819
3 6 77 0 0 12416 0 80 85 0 0 4
368 331
537 331
537 717
995 717
3 6 78 0 0 12416 0 81 86 0 0 4
317 295
550 295
550 617
995 617
1 2 21 0 0 0 0 96 64 0 0 3
61 66
61 778
111 778
2 1 24 0 0 0 0 96 64 0 0 3
55 66
55 760
111 760
2 2 24 0 0 0 0 65 96 0 0 3
113 728
55 728
55 66
3 1 23 0 0 0 0 96 65 0 0 3
49 66
49 710
113 710
3 2 23 0 0 0 0 96 66 0 0 3
49 66
49 676
111 676
4 1 31 0 0 0 0 96 66 0 0 3
43 66
43 658
111 658
3 8 79 0 0 4224 0 67 87 0 0 4
159 612
605 612
605 528
995 528
4 2 31 0 0 0 0 96 67 0 0 3
43 66
43 621
110 621
1 1 80 0 0 4224 0 93 67 0 0 3
24 64
24 603
110 603
3 8 81 0 0 4224 0 68 88 0 0 4
166 564
599 564
599 425
996 425
3 8 82 0 0 4224 0 69 89 0 0 4
159 513
592 513
592 323
1002 323
3 8 83 0 0 12416 0 70 90 0 0 4
233 448
583 448
583 223
1001 223
2 1 80 0 0 0 0 68 93 0 0 3
117 573
24 573
24 64
2 1 84 0 0 4224 0 93 68 0 0 3
18 64
18 555
117 555
2 2 84 0 0 0 0 69 93 0 0 3
110 522
18 522
18 64
3 1 85 0 0 4224 0 93 69 0 0 3
12 64
12 504
110 504
2 3 85 0 0 0 0 70 93 0 0 3
184 457
12 457
12 64
3 6 86 0 0 12416 0 82 87 0 0 4
270 266
518 266
518 510
995 510
3 6 87 0 0 12416 0 83 88 0 0 4
219 225
501 225
501 407
996 407
3 6 88 0 0 12416 0 95 89 0 0 4
171 193
511 193
511 305
1002 305
3 6 89 0 0 12416 0 94 90 0 0 4
122 163
516 163
516 205
1001 205
4 8 72 0 0 8320 0 93 92 0 0 3
6 64
6 130
1001 130
4 6 72 0 0 0 0 93 92 0 0 3
6 64
6 112
1001 112
14 1 90 0 0 8320 0 84 71 0 0 3
1055 837
1417 837
1417 52
14 1 11 0 0 8320 0 85 72 0 0 3
1059 735
1382 735
1382 42
14 1 12 0 0 8320 0 86 73 0 0 3
1059 635
1354 635
1354 41
14 1 13 0 0 0 0 87 74 0 0 3
1059 528
1332 528
1332 41
14 1 14 0 0 0 0 88 75 0 0 3
1060 425
1298 425
1298 45
14 1 16 0 0 0 0 89 76 0 0 3
1066 323
1273 323
1273 49
14 1 17 0 0 0 0 90 77 0 0 3
1065 223
1250 223
1250 51
14 1 18 0 0 0 0 92 78 0 0 3
1065 130
1215 130
1215 52
2 1 21 0 0 0 0 79 96 0 0 3
369 364
61 364
61 66
3 1 77 0 0 0 0 80 79 0 0 4
368 331
366 331
366 346
369 346
2 2 24 0 0 0 0 80 96 0 0 3
319 340
55 340
55 66
3 1 78 0 0 0 0 81 80 0 0 3
317 295
317 322
319 322
2 3 23 0 0 0 0 81 96 0 0 3
268 304
49 304
49 66
3 1 86 0 0 0 0 82 81 0 0 3
270 266
268 266
268 286
4 2 31 0 0 0 0 96 82 0 0 3
43 66
43 275
221 275
3 1 87 0 0 0 0 83 82 0 0 4
219 225
220 225
220 257
221 257
1 2 80 0 0 0 0 93 83 0 0 3
24 64
24 234
170 234
3 1 88 0 0 0 0 95 83 0 0 4
171 193
169 193
169 216
170 216
2 2 84 0 0 0 0 93 95 0 0 3
18 64
18 202
122 202
12 1 91 0 0 8320 0 84 3 0 0 3
1061 801
1160 801
1160 34
12 1 91 0 0 0 0 85 3 0 0 3
1065 699
1160 699
1160 34
12 1 91 0 0 0 0 86 3 0 0 3
1065 599
1160 599
1160 34
12 1 91 0 0 0 0 87 3 0 0 3
1065 492
1160 492
1160 34
12 1 91 0 0 0 0 88 3 0 0 3
1066 389
1160 389
1160 34
12 1 91 0 0 0 0 89 3 0 0 3
1072 287
1160 287
1160 34
12 1 91 0 0 0 0 90 3 0 0 3
1071 187
1160 187
1160 34
1 12 91 0 0 0 0 3 92 0 0 3
1160 34
1160 94
1071 94
9 3 92 0 0 8192 0 86 91 0 0 3
1059 572
1112 572
1112 57
9 3 92 0 0 8192 0 85 91 0 0 3
1059 672
1112 672
1112 57
3 9 92 0 0 4224 0 91 84 0 0 3
1112 57
1112 774
1055 774
10 2 93 0 0 8320 0 84 91 0 0 3
1055 783
1118 783
1118 57
10 2 93 0 0 0 0 85 91 0 0 3
1059 681
1118 681
1118 57
2 10 93 0 0 0 0 91 86 0 0 3
1118 57
1118 581
1059 581
11 1 94 0 0 8320 0 84 91 0 0 3
1055 792
1124 792
1124 57
11 1 94 0 0 0 0 85 91 0 0 3
1059 690
1124 690
1124 57
11 1 94 0 0 0 0 86 91 0 0 3
1059 590
1124 590
1124 57
9 3 92 0 0 0 0 87 91 0 0 3
1059 465
1112 465
1112 57
9 3 92 0 0 0 0 88 91 0 0 3
1060 362
1112 362
1112 57
2 10 93 0 0 0 0 91 87 0 0 3
1118 57
1118 474
1059 474
2 10 93 0 0 0 0 91 88 0 0 3
1118 57
1118 371
1060 371
11 1 94 0 0 0 0 87 91 0 0 3
1059 483
1124 483
1124 57
1 11 94 0 0 0 0 91 88 0 0 3
1124 57
1124 380
1060 380
1 11 94 0 0 0 0 91 89 0 0 3
1124 57
1124 278
1066 278
10 2 93 0 0 0 0 89 91 0 0 3
1066 269
1118 269
1118 57
3 9 92 0 0 0 0 91 89 0 0 3
1112 57
1112 260
1066 260
11 1 94 0 0 0 0 90 91 0 0 3
1065 178
1124 178
1124 57
2 10 93 0 0 0 0 91 90 0 0 3
1118 57
1118 169
1065 169
9 3 92 0 0 0 0 90 91 0 0 3
1065 160
1112 160
1112 57
3 9 92 0 0 0 0 91 92 0 0 3
1112 57
1112 67
1065 67
2 10 93 0 0 0 0 91 92 0 0 3
1118 57
1118 76
1065 76
1 11 94 0 0 0 0 91 92 0 0 3
1124 57
1124 85
1065 85
3 1 85 0 0 0 0 93 94 0 0 3
12 64
12 154
73 154
4 2 72 0 0 0 0 93 94 0 0 3
6 64
6 172
73 172
3 1 89 0 0 0 0 94 95 0 0 2
122 163
122 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
