CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 600 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
50
13 Logic Switch~
5 789 992 0 1 11
0 19
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45437.7 0
0
13 Logic Switch~
5 1160 22 0 1 11
0 45
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
45437.7 1
0
9 Inverter~
13 102 1075 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3124 0 0
2
45437.8 0
0
9 Inverter~
13 113 1046 0 2 22
0 7 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3421 0 0
2
45437.8 0
0
9 Inverter~
13 157 1037 0 2 22
0 8 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
8157 0 0
2
45437.8 0
0
9 Inverter~
13 118 979 0 2 22
0 4 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
5572 0 0
2
45437.8 0
0
9 Inverter~
13 92 928 0 2 22
0 12 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
8901 0 0
2
45437.8 0
0
9 Inverter~
13 157 946 0 2 22
0 7 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
7361 0 0
2
45437.8 0
0
7 Ground~
168 990 922 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4747 0 0
2
45437.8 0
0
5 7415~
219 381 1084 0 4 22
0 3 8 12 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U17B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 12 0
1 U
972 0 0
2
45437.8 0
0
5 7415~
219 381 1037 0 4 22
0 4 6 5 16
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U17A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 12 0
1 U
3472 0 0
2
45437.8 0
0
9 2-In AND~
219 378 937 0 3 22
0 11 10 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
9998 0 0
2
45437.8 0
0
9 2-In AND~
219 380 988 0 3 22
0 9 7 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3536 0 0
2
45437.8 0
0
8 4-In OR~
219 573 902 0 5 22
0 18 17 16 15 14
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
4597 0 0
2
45437.8 0
0
9 CC 7-Seg~
183 833 926 0 16 19
10 14 49 50 51 52 53 54 19 2
1 2 2 2 2 2 2
0
0 0 21104 270
5 REDCC
16 -41 51 -33
5 DISP3
-21 -39 14 -31
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3835 0 0
2
45437.7 0
0
6 74136~
219 127 769 0 3 22
0 7 12 20
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3670 0 0
2
45437.7 0
0
6 74136~
219 129 719 0 3 22
0 8 7 21
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5616 0 0
2
45437.7 0
0
6 74136~
219 127 667 0 3 22
0 4 8 22
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
9323 0 0
2
45437.7 0
0
6 74136~
219 126 612 0 3 22
0 27 4 26
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
317 0 0
2
45437.7 0
0
6 74136~
219 133 564 0 3 22
0 31 27 28
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3108 0 0
2
45437.7 0
0
6 74136~
219 126 513 0 3 22
0 32 31 29
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4299 0 0
2
45437.7 0
0
6 74136~
219 200 448 0 3 22
0 13 32 30
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9672 0 0
2
45437.7 0
0
14 Logic Display~
6 1417 34 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90125e-315 0
0
14 Logic Display~
6 1382 24 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.90125e-315 5.26354e-315
0
14 Logic Display~
6 1354 23 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.90125e-315 5.30499e-315
0
14 Logic Display~
6 1332 23 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.90125e-315 5.32571e-315
0
14 Logic Display~
6 1298 27 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90125e-315 5.34643e-315
0
14 Logic Display~
6 1273 31 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90125e-315 5.3568e-315
0
14 Logic Display~
6 1250 33 0 1 2
10 43
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90125e-315 5.36716e-315
0
14 Logic Display~
6 1215 34 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.90125e-315 5.37752e-315
0
6 74136~
219 385 355 0 3 22
0 24 12 23
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3409 0 0
2
5.90125e-315 5.38788e-315
0
6 74136~
219 335 331 0 3 22
0 25 7 24
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3951 0 0
2
5.90125e-315 5.39306e-315
0
6 74136~
219 284 295 0 3 22
0 33 8 25
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8885 0 0
2
5.90125e-315 5.39824e-315
0
6 74136~
219 237 266 0 3 22
0 34 4 33
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3780 0 0
2
5.90125e-315 5.40342e-315
0
6 74136~
219 186 225 0 3 22
0 35 27 34
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9265 0 0
2
5.90125e-315 5.4086e-315
0
7 74LS251
144 1023 801 0 14 29
0 55 56 57 58 59 23 60 20 46
47 48 45 61 37
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9442 0 0
2
45437.7 4
0
7 74LS251
144 1027 699 0 14 29
0 62 63 64 65 66 24 67 21 46
47 48 45 68 38
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9424 0 0
2
45437.7 5
0
7 74LS251
144 1027 599 0 14 29
0 69 70 71 72 73 25 74 22 46
47 48 45 75 39
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9968 0 0
2
45437.7 6
0
7 74LS251
144 1027 492 0 14 29
0 76 77 78 79 80 33 81 26 46
47 48 45 82 40
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9281 0 0
2
45437.7 7
0
7 74LS251
144 1028 389 0 14 29
0 83 84 85 86 87 34 88 28 46
47 48 45 89 41
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8464 0 0
2
45437.7 8
0
7 74LS251
144 1034 287 0 14 29
0 90 91 92 93 94 35 95 29 46
47 48 45 96 42
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7168 0 0
2
45437.7 9
0
7 74LS251
144 1033 187 0 14 29
0 97 98 99 100 101 36 102 30 46
47 48 45 103 43
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3171 0 0
2
45437.7 10
0
8 Hex Key~
166 1115 33 0 11 12
0 48 47 46 104 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
4139 0 0
2
45437.7 11
0
7 74LS251
144 1033 94 0 14 29
0 105 106 107 108 109 13 110 13 46
47 48 45 111 44
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6435 0 0
2
45437.7 12
0
12 Hex Display~
7 1859 45 0 18 19
10 37 38 39 40 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5283 0 0
2
45437.7 13
0
8 Hex Key~
166 15 40 0 11 12
0 27 31 32 13 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6874 0 0
2
45437.7 14
0
6 74136~
219 89 163 0 3 22
0 32 13 36
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5305 0 0
2
45437.7 15
0
12 Hex Display~
7 1799 42 0 18 19
10 41 42 43 44 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
34 0 0
2
45437.7 16
0
6 74136~
219 138 193 0 3 22
0 36 31 35
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
969 0 0
2
45437.7 17
0
8 Hex Key~
166 52 42 0 11 12
0 12 7 8 4 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8402 0 0
2
45437.7 18
0
115
1 9 0 0 0 0 0 9 15 0 0 2
983 923
872 923
1 5 0 0 0 0 0 15 14 0 0 2
794 902
606 902
8 1 0 0 0 0 0 15 1 0 0 3
794 944
790 944
790 979
2 1 3 0 0 12416 0 3 10 0 0 2
123 1075
357 1075
4 1 4 0 0 4224 0 50 3 0 0 3
43 66
43 1075
87 1075
3 2 5 0 0 4224 0 11 4 0 0 2
357 1046
134 1046
2 2 6 0 0 4224 0 5 11 0 0 2
178 1037
357 1037
2 1 7 0 0 4224 0 50 4 0 0 3
55 66
55 1046
98 1046
3 1 8 0 0 4096 0 50 5 0 0 3
49 66
49 1037
142 1037
2 2 7 0 0 0 0 50 13 0 0 3
55 66
55 997
356 997
2 1 9 0 0 4224 0 6 13 0 0 2
139 979
356 979
4 1 4 0 0 0 0 50 6 0 0 3
43 66
43 979
103 979
2 2 10 0 0 4224 0 12 8 0 0 2
354 946
178 946
2 1 11 0 0 4224 0 7 12 0 0 2
113 928
354 928
1 1 12 0 0 4096 0 50 7 0 0 3
61 66
61 928
77 928
2 1 7 0 0 0 0 50 8 0 0 3
55 66
55 946
142 946
4 1 13 0 0 4096 0 46 22 0 0 3
6 64
6 439
184 439
4 4 15 0 0 12416 0 14 10 0 0 4
556 916
536 916
536 1084
402 1084
4 3 16 0 0 8320 0 11 14 0 0 4
402 1037
512 1037
512 907
556 907
2 3 17 0 0 8320 0 14 13 0 0 4
556 898
474 898
474 988
401 988
3 1 18 0 0 12432 0 12 14 0 0 4
399 937
457 937
457 889
556 889
1 3 12 0 0 4224 0 50 10 0 0 3
61 66
61 1093
357 1093
2 3 8 0 0 8320 0 10 50 0 0 3
357 1084
49 1084
49 66
4 1 4 0 0 0 0 50 11 0 0 3
43 66
43 1028
357 1028
3 8 20 0 0 4224 0 16 36 0 0 4
160 769
603 769
603 837
991 837
3 8 21 0 0 16512 0 17 37 0 0 5
162 719
162 724
577 724
577 735
995 735
3 8 22 0 0 12416 0 18 38 0 0 4
160 667
566 667
566 635
995 635
3 6 23 0 0 8320 0 31 36 0 0 4
418 355
528 355
528 819
991 819
3 6 24 0 0 12416 0 32 37 0 0 4
368 331
537 331
537 717
995 717
3 6 25 0 0 12416 0 33 38 0 0 4
317 295
550 295
550 617
995 617
1 2 12 0 0 128 0 50 16 0 0 3
61 66
61 778
111 778
2 1 7 0 0 128 0 50 16 0 0 3
55 66
55 760
111 760
2 2 7 0 0 0 0 17 50 0 0 3
113 728
55 728
55 66
3 1 8 0 0 128 0 50 17 0 0 3
49 66
49 710
113 710
3 2 8 0 0 0 0 50 18 0 0 3
49 66
49 676
111 676
4 1 4 0 0 128 0 50 18 0 0 3
43 66
43 658
111 658
3 8 26 0 0 4224 0 19 39 0 0 4
159 612
605 612
605 528
995 528
4 2 4 0 0 0 0 50 19 0 0 3
43 66
43 621
110 621
1 1 27 0 0 4224 0 46 19 0 0 3
24 64
24 603
110 603
3 8 28 0 0 4224 0 20 40 0 0 4
166 564
599 564
599 425
996 425
3 8 29 0 0 4224 0 21 41 0 0 4
159 513
592 513
592 323
1002 323
3 8 30 0 0 12416 0 22 42 0 0 4
233 448
583 448
583 223
1001 223
2 1 27 0 0 0 0 20 46 0 0 3
117 573
24 573
24 64
2 1 31 0 0 4224 0 46 20 0 0 3
18 64
18 555
117 555
2 2 31 0 0 0 0 21 46 0 0 3
110 522
18 522
18 64
3 1 32 0 0 4224 0 46 21 0 0 3
12 64
12 504
110 504
2 3 32 0 0 0 0 22 46 0 0 3
184 457
12 457
12 64
3 6 33 0 0 12416 0 34 39 0 0 4
270 266
518 266
518 510
995 510
3 6 34 0 0 12416 0 35 40 0 0 4
219 225
501 225
501 407
996 407
3 6 35 0 0 12416 0 49 41 0 0 4
171 193
511 193
511 305
1002 305
3 6 36 0 0 12416 0 47 42 0 0 4
122 163
516 163
516 205
1001 205
4 8 13 0 0 8320 0 46 44 0 0 3
6 64
6 130
1001 130
4 6 13 0 0 0 0 46 44 0 0 3
6 64
6 112
1001 112
14 1 37 0 0 8192 0 36 23 0 0 3
1055 837
1417 837
1417 52
14 1 38 0 0 8192 0 37 24 0 0 3
1059 735
1382 735
1382 42
14 1 39 0 0 8192 0 38 25 0 0 3
1059 635
1354 635
1354 41
14 1 40 0 0 8192 0 39 26 0 0 3
1059 528
1332 528
1332 41
14 1 41 0 0 8192 0 40 27 0 0 3
1060 425
1298 425
1298 45
14 1 42 0 0 8192 0 41 28 0 0 3
1066 323
1273 323
1273 49
14 1 43 0 0 4096 0 42 29 0 0 3
1065 223
1250 223
1250 51
14 1 44 0 0 4096 0 44 30 0 0 3
1065 130
1215 130
1215 52
14 1 37 0 0 4224 0 36 45 0 0 3
1055 837
1868 837
1868 69
14 2 38 0 0 4224 0 37 45 0 0 3
1059 735
1862 735
1862 69
14 3 39 0 0 4224 0 38 45 0 0 3
1059 635
1856 635
1856 69
14 4 40 0 0 4224 0 39 45 0 0 3
1059 528
1850 528
1850 69
2 1 12 0 0 128 0 31 50 0 0 3
369 364
61 364
61 66
3 1 24 0 0 0 0 32 31 0 0 4
368 331
366 331
366 346
369 346
2 2 7 0 0 128 0 32 50 0 0 3
319 340
55 340
55 66
3 1 25 0 0 0 0 33 32 0 0 3
317 295
317 322
319 322
2 3 8 0 0 128 0 33 50 0 0 3
268 304
49 304
49 66
3 1 33 0 0 0 0 34 33 0 0 3
270 266
268 266
268 286
4 2 4 0 0 128 0 50 34 0 0 3
43 66
43 275
221 275
3 1 34 0 0 0 0 35 34 0 0 4
219 225
220 225
220 257
221 257
1 2 27 0 0 128 0 46 35 0 0 3
24 64
24 234
170 234
3 1 35 0 0 0 0 49 35 0 0 4
171 193
169 193
169 216
170 216
2 2 31 0 0 128 0 46 49 0 0 3
18 64
18 202
122 202
12 1 45 0 0 8320 0 36 2 0 0 3
1061 801
1160 801
1160 34
12 1 45 0 0 0 0 37 2 0 0 3
1065 699
1160 699
1160 34
12 1 45 0 0 0 0 38 2 0 0 3
1065 599
1160 599
1160 34
12 1 45 0 0 0 0 39 2 0 0 3
1065 492
1160 492
1160 34
12 1 45 0 0 0 0 40 2 0 0 3
1066 389
1160 389
1160 34
12 1 45 0 0 0 0 41 2 0 0 3
1072 287
1160 287
1160 34
12 1 45 0 0 0 0 42 2 0 0 3
1071 187
1160 187
1160 34
1 12 45 0 0 0 0 2 44 0 0 3
1160 34
1160 94
1071 94
14 1 41 0 0 4224 0 40 48 0 0 3
1060 425
1808 425
1808 66
14 2 42 0 0 4224 0 41 48 0 0 3
1066 323
1802 323
1802 66
14 3 43 0 0 4224 0 42 48 0 0 3
1065 223
1796 223
1796 66
14 4 44 0 0 4224 0 44 48 0 0 3
1065 130
1790 130
1790 66
9 3 46 0 0 8192 0 38 43 0 0 3
1059 572
1112 572
1112 57
9 3 46 0 0 8192 0 37 43 0 0 3
1059 672
1112 672
1112 57
3 9 46 0 0 4224 0 43 36 0 0 3
1112 57
1112 774
1055 774
10 2 47 0 0 8320 0 36 43 0 0 3
1055 783
1118 783
1118 57
10 2 47 0 0 0 0 37 43 0 0 3
1059 681
1118 681
1118 57
2 10 47 0 0 0 0 43 38 0 0 3
1118 57
1118 581
1059 581
11 1 48 0 0 8320 0 36 43 0 0 3
1055 792
1124 792
1124 57
11 1 48 0 0 0 0 37 43 0 0 3
1059 690
1124 690
1124 57
11 1 48 0 0 0 0 38 43 0 0 3
1059 590
1124 590
1124 57
9 3 46 0 0 0 0 39 43 0 0 3
1059 465
1112 465
1112 57
9 3 46 0 0 0 0 40 43 0 0 3
1060 362
1112 362
1112 57
2 10 47 0 0 0 0 43 39 0 0 3
1118 57
1118 474
1059 474
2 10 47 0 0 0 0 43 40 0 0 3
1118 57
1118 371
1060 371
11 1 48 0 0 0 0 39 43 0 0 3
1059 483
1124 483
1124 57
1 11 48 0 0 0 0 43 40 0 0 3
1124 57
1124 380
1060 380
1 11 48 0 0 0 0 43 41 0 0 3
1124 57
1124 278
1066 278
10 2 47 0 0 0 0 41 43 0 0 3
1066 269
1118 269
1118 57
3 9 46 0 0 0 0 43 41 0 0 3
1112 57
1112 260
1066 260
11 1 48 0 0 0 0 42 43 0 0 3
1065 178
1124 178
1124 57
2 10 47 0 0 0 0 43 42 0 0 3
1118 57
1118 169
1065 169
9 3 46 0 0 0 0 42 43 0 0 3
1065 160
1112 160
1112 57
3 9 46 0 0 0 0 43 44 0 0 3
1112 57
1112 67
1065 67
2 10 47 0 0 0 0 43 44 0 0 3
1118 57
1118 76
1065 76
1 11 48 0 0 0 0 43 44 0 0 3
1124 57
1124 85
1065 85
3 1 32 0 0 128 0 46 47 0 0 3
12 64
12 154
73 154
4 2 13 0 0 0 0 46 47 0 0 3
6 64
6 172
73 172
3 1 36 0 0 0 0 47 49 0 0 2
122 163
122 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
