CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
500 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 1160 22 0 1 11
0 33
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90124e-315 0
0
6 74136~
219 140 715 0 3 22
0 6 5 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
391 0 0
2
45435.5 0
0
6 74136~
219 134 671 0 3 22
0 7 6 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3124 0 0
2
45435.5 0
0
6 74136~
219 137 623 0 3 22
0 9 7 8
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3421 0 0
2
45435.5 0
0
6 74136~
219 138 565 0 3 22
0 10 9 11
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
8157 0 0
2
45435.5 0
0
6 74136~
219 140 516 0 3 22
0 16 10 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
5572 0 0
2
45435.5 0
0
6 74136~
219 138 469 0 3 22
0 17 17 13
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8901 0 0
2
45435.5 0
0
6 74136~
219 136 417 0 3 22
0 15 17 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7361 0 0
2
45435.5 0
0
7 Ground~
168 1525 9 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.90124e-315 0
0
9 CC 7-Seg~
183 1536 77 0 17 19
10 37 38 39 40 41 42 43 44 2
2 2 2 2 2 2 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1417 34 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
45435.5 0
0
14 Logic Display~
6 1382 24 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
45435.5 1
0
14 Logic Display~
6 1354 23 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
45435.5 2
0
14 Logic Display~
6 1332 23 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
45435.5 3
0
14 Logic Display~
6 1298 27 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
45435.5 4
0
14 Logic Display~
6 1273 31 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
45435.5 5
0
14 Logic Display~
6 1250 33 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
45435.5 6
0
14 Logic Display~
6 1215 34 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
45435.5 7
0
6 74136~
219 385 355 0 3 22
0 19 5 18
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
317 0 0
2
45435.5 8
0
6 74136~
219 335 331 0 3 22
0 20 6 19
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3108 0 0
2
45435.5 9
0
6 74136~
219 284 295 0 3 22
0 21 7 20
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
45435.5 10
0
6 74136~
219 237 266 0 3 22
0 22 9 21
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
45435.5 11
0
6 74136~
219 186 225 0 3 22
0 23 10 22
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7876 0 0
2
45435.5 12
0
12 Hex Display~
7 585 27 0 18 19
10 18 19 20 21 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6369 0 0
2
45435.5 13
0
12 Hex Display~
7 533 28 0 18 19
10 22 23 24 15 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9172 0 0
2
45435.5 14
0
7 74LS251
144 1023 801 0 14 29
0 45 46 47 48 49 18 50 3 34
35 36 33 51 25
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
5.90124e-315 5.26354e-315
0
7 74LS251
144 1027 699 0 14 29
0 52 53 54 55 56 19 57 4 34
35 36 33 58 26
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3820 0 0
2
5.90124e-315 5.30499e-315
0
7 74LS251
144 1027 599 0 14 29
0 59 60 61 62 63 20 64 8 34
35 36 33 65 27
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7678 0 0
2
5.90124e-315 5.32571e-315
0
7 74LS251
144 1027 492 0 14 29
0 66 67 68 69 70 21 71 11 34
35 36 33 72 28
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
961 0 0
2
5.90124e-315 5.34643e-315
0
7 74LS251
144 1028 389 0 14 29
0 73 74 75 76 77 22 78 12 34
35 36 33 79 29
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3178 0 0
2
5.90124e-315 5.3568e-315
0
7 74LS251
144 1034 287 0 14 29
0 80 81 82 83 84 23 85 13 34
35 36 33 86 30
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
5.90124e-315 5.36716e-315
0
7 74LS251
144 1033 187 0 14 29
0 87 88 89 90 91 24 92 14 34
35 36 33 93 31
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3951 0 0
2
5.90124e-315 5.37752e-315
0
8 Hex Key~
166 1115 33 0 11 12
0 36 35 34 94 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8885 0 0
2
5.90124e-315 5.38788e-315
0
7 74LS251
144 1033 94 0 14 29
0 95 96 97 98 99 15 100 15 34
35 36 33 101 32
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3780 0 0
2
5.90124e-315 5.39306e-315
0
12 Hex Display~
7 1859 45 0 16 19
10 25 26 27 28 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9265 0 0
2
5.90124e-315 5.39824e-315
0
8 Hex Key~
166 15 40 0 11 12
0 10 16 17 15 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9442 0 0
2
5.90124e-315 5.40342e-315
0
6 74136~
219 89 163 0 3 22
0 17 15 24
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9424 0 0
2
5.90124e-315 5.4086e-315
0
12 Hex Display~
7 1799 42 0 18 19
10 29 30 31 32 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9968 0 0
2
5.90124e-315 5.41378e-315
0
6 74136~
219 138 193 0 3 22
0 24 16 23
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9281 0 0
2
5.90124e-315 5.41896e-315
0
8 Hex Key~
166 52 42 0 11 12
0 5 6 7 9 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8464 0 0
2
5.90124e-315 5.42414e-315
0
101
3 8 3 0 0 12416 0 2 26 0 0 4
173 715
181 715
181 837
991 837
3 8 4 0 0 12432 0 3 27 0 0 4
167 671
203 671
203 735
995 735
1 2 5 0 0 4224 0 40 2 0 0 3
61 66
61 724
124 724
2 1 6 0 0 4224 0 40 2 0 0 3
55 66
55 706
124 706
2 2 6 0 0 0 0 40 3 0 0 3
55 66
55 680
118 680
3 1 7 0 0 4224 0 40 3 0 0 3
49 66
49 662
118 662
3 8 8 0 0 12416 0 4 28 0 0 4
170 623
180 623
180 635
995 635
3 2 7 0 0 0 0 40 4 0 0 3
49 66
49 632
121 632
4 1 9 0 0 4224 0 40 4 0 0 3
43 66
43 614
121 614
4 2 9 0 0 0 0 40 5 0 0 3
43 66
43 574
122 574
1 1 10 0 0 8320 0 5 36 0 0 3
122 556
24 556
24 64
3 8 11 0 0 4224 0 5 29 0 0 4
171 565
987 565
987 528
995 528
3 8 12 0 0 8320 0 6 30 0 0 3
173 516
173 425
996 425
3 8 13 0 0 4224 0 7 31 0 0 4
171 469
652 469
652 323
1002 323
3 8 14 0 0 8320 0 8 32 0 0 5
169 417
169 392
625 392
625 223
1001 223
4 8 15 0 0 8320 0 36 34 0 0 3
6 64
6 130
1001 130
1 2 10 0 0 0 0 36 6 0 0 3
24 64
24 525
124 525
2 1 16 0 0 4224 0 36 6 0 0 3
18 64
18 507
124 507
3 2 17 0 0 4224 0 36 7 0 0 3
12 64
12 478
122 478
3 1 17 0 0 0 0 36 7 0 0 3
12 64
12 460
122 460
3 2 17 0 0 0 0 36 8 0 0 3
12 64
12 426
120 426
4 1 15 0 0 0 0 36 8 0 0 3
6 64
6 408
120 408
9 1 2 0 0 8320 0 10 9 0 0 4
1536 35
1536 25
1525 25
1525 17
3 6 18 0 0 8320 0 19 26 0 0 4
418 355
594 355
594 819
991 819
3 6 19 0 0 12416 0 20 27 0 0 4
368 331
588 331
588 717
995 717
3 6 20 0 0 12416 0 21 28 0 0 4
317 295
582 295
582 617
995 617
3 6 21 0 0 12416 0 22 29 0 0 4
270 266
576 266
576 510
995 510
3 6 22 0 0 12416 0 23 30 0 0 4
219 225
603 225
603 407
996 407
3 6 23 0 0 4224 0 39 31 0 0 4
171 193
652 193
652 305
1002 305
3 6 24 0 0 4224 0 37 32 0 0 4
122 163
678 163
678 205
1001 205
4 6 15 0 0 128 0 36 34 0 0 3
6 64
6 112
1001 112
14 1 25 0 0 8192 0 26 11 0 0 3
1055 837
1417 837
1417 52
14 1 26 0 0 8192 0 27 12 0 0 3
1059 735
1382 735
1382 42
14 1 27 0 0 8192 0 28 13 0 0 3
1059 635
1354 635
1354 41
14 1 28 0 0 8192 0 29 14 0 0 3
1059 528
1332 528
1332 41
14 1 29 0 0 8192 0 30 15 0 0 3
1060 425
1298 425
1298 45
14 1 30 0 0 8192 0 31 16 0 0 3
1066 323
1273 323
1273 49
14 1 31 0 0 4096 0 32 17 0 0 3
1065 223
1250 223
1250 51
14 1 32 0 0 4096 0 34 18 0 0 3
1065 130
1215 130
1215 52
14 1 25 0 0 4224 0 26 35 0 0 3
1055 837
1868 837
1868 69
14 2 26 0 0 4224 0 27 35 0 0 3
1059 735
1862 735
1862 69
14 3 27 0 0 4224 0 28 35 0 0 3
1059 635
1856 635
1856 69
14 4 28 0 0 4224 0 29 35 0 0 3
1059 528
1850 528
1850 69
3 1 18 0 0 0 0 19 24 0 0 3
418 355
594 355
594 51
2 1 5 0 0 128 0 19 40 0 0 3
369 364
61 364
61 66
3 1 19 0 0 0 0 20 19 0 0 4
368 331
366 331
366 346
369 346
3 2 19 0 0 0 0 20 24 0 0 3
368 331
588 331
588 51
2 2 6 0 0 128 0 20 40 0 0 3
319 340
55 340
55 66
3 1 20 0 0 0 0 21 20 0 0 3
317 295
317 322
319 322
3 3 20 0 0 0 0 21 24 0 0 3
317 295
582 295
582 51
2 3 7 0 0 128 0 21 40 0 0 3
268 304
49 304
49 66
3 1 21 0 0 0 0 22 21 0 0 3
270 266
268 266
268 286
3 4 21 0 0 0 0 22 24 0 0 3
270 266
576 266
576 51
4 2 9 0 0 128 0 40 22 0 0 3
43 66
43 275
221 275
3 1 22 0 0 0 0 23 22 0 0 4
219 225
220 225
220 257
221 257
3 1 22 0 0 0 0 23 25 0 0 3
219 225
542 225
542 52
1 2 10 0 0 128 0 36 23 0 0 3
24 64
24 234
170 234
3 1 23 0 0 0 0 39 23 0 0 4
171 193
169 193
169 216
170 216
3 2 23 0 0 0 0 39 25 0 0 3
171 193
536 193
536 52
2 2 16 0 0 128 0 36 39 0 0 3
18 64
18 202
122 202
3 3 24 0 0 0 0 37 25 0 0 3
122 163
530 163
530 52
4 4 15 0 0 0 0 36 25 0 0 4
6 64
6 130
524 130
524 52
12 1 33 0 0 8320 0 26 1 0 0 3
1061 801
1160 801
1160 34
12 1 33 0 0 0 0 27 1 0 0 3
1065 699
1160 699
1160 34
12 1 33 0 0 0 0 28 1 0 0 3
1065 599
1160 599
1160 34
12 1 33 0 0 0 0 29 1 0 0 3
1065 492
1160 492
1160 34
12 1 33 0 0 0 0 30 1 0 0 3
1066 389
1160 389
1160 34
12 1 33 0 0 0 0 31 1 0 0 3
1072 287
1160 287
1160 34
12 1 33 0 0 0 0 32 1 0 0 3
1071 187
1160 187
1160 34
1 12 33 0 0 0 0 1 34 0 0 3
1160 34
1160 94
1071 94
14 1 29 0 0 4224 0 30 38 0 0 3
1060 425
1808 425
1808 66
14 2 30 0 0 4224 0 31 38 0 0 3
1066 323
1802 323
1802 66
14 3 31 0 0 4224 0 32 38 0 0 3
1065 223
1796 223
1796 66
14 4 32 0 0 4224 0 34 38 0 0 3
1065 130
1790 130
1790 66
9 3 34 0 0 8192 0 28 33 0 0 3
1059 572
1112 572
1112 57
9 3 34 0 0 8192 0 27 33 0 0 3
1059 672
1112 672
1112 57
3 9 34 0 0 4224 0 33 26 0 0 3
1112 57
1112 774
1055 774
10 2 35 0 0 8320 0 26 33 0 0 3
1055 783
1118 783
1118 57
10 2 35 0 0 0 0 27 33 0 0 3
1059 681
1118 681
1118 57
2 10 35 0 0 0 0 33 28 0 0 3
1118 57
1118 581
1059 581
11 1 36 0 0 8320 0 26 33 0 0 3
1055 792
1124 792
1124 57
11 1 36 0 0 0 0 27 33 0 0 3
1059 690
1124 690
1124 57
11 1 36 0 0 0 0 28 33 0 0 3
1059 590
1124 590
1124 57
9 3 34 0 0 0 0 29 33 0 0 3
1059 465
1112 465
1112 57
9 3 34 0 0 0 0 30 33 0 0 3
1060 362
1112 362
1112 57
2 10 35 0 0 0 0 33 29 0 0 3
1118 57
1118 474
1059 474
2 10 35 0 0 0 0 33 30 0 0 3
1118 57
1118 371
1060 371
11 1 36 0 0 0 0 29 33 0 0 3
1059 483
1124 483
1124 57
1 11 36 0 0 0 0 33 30 0 0 3
1124 57
1124 380
1060 380
1 11 36 0 0 0 0 33 31 0 0 3
1124 57
1124 278
1066 278
10 2 35 0 0 0 0 31 33 0 0 3
1066 269
1118 269
1118 57
3 9 34 0 0 0 0 33 31 0 0 3
1112 57
1112 260
1066 260
11 1 36 0 0 0 0 32 33 0 0 3
1065 178
1124 178
1124 57
2 10 35 0 0 0 0 33 32 0 0 3
1118 57
1118 169
1065 169
9 3 34 0 0 0 0 32 33 0 0 3
1065 160
1112 160
1112 57
3 9 34 0 0 0 0 33 34 0 0 3
1112 57
1112 67
1065 67
2 10 35 0 0 0 0 33 34 0 0 3
1118 57
1118 76
1065 76
1 11 36 0 0 0 0 33 34 0 0 3
1124 57
1124 85
1065 85
3 1 17 0 0 128 0 36 37 0 0 3
12 64
12 154
73 154
4 2 15 0 0 0 0 36 37 0 0 3
6 64
6 172
73 172
3 1 24 0 0 0 0 37 39 0 0 2
122 163
122 184
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
152 429 243 453
164 438 230 454
11 Codificador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
223 192 330 216
234 201 318 217
14 DE_Codificador
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
