CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 427 589 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
45435.4 0
0
13 Logic Switch~
5 1160 22 0 1 11
0 26
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9442 0 0
2
45435.4 0
0
7 Ground~
168 482 380 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9424 0 0
2
45435.4 0
0
9 CC 7-Seg~
183 482 491 0 17 19
10 31 32 33 34 35 3 36 37 2
2 2 2 2 2 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9968 0 0
2
45435.4 0
0
14 Logic Display~
6 1417 34 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1382 24 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1354 23 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1332 23 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1298 27 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1273 31 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1250 33 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 1215 34 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.90124e-315 0
0
6 74136~
219 385 355 0 3 22
0 14 19 13
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5305 0 0
2
5.90124e-315 0
0
6 74136~
219 335 331 0 3 22
0 15 20 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
34 0 0
2
5.90124e-315 0
0
6 74136~
219 284 295 0 3 22
0 16 21 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
969 0 0
2
5.90124e-315 0
0
6 74136~
219 237 266 0 3 22
0 17 22 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8402 0 0
2
5.90124e-315 0
0
6 74136~
219 186 225 0 3 22
0 18 23 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3751 0 0
2
5.90124e-315 0
0
12 Hex Display~
7 585 27 0 18 19
10 13 14 15 16 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4292 0 0
2
5.90124e-315 0
0
12 Hex Display~
7 533 28 0 18 19
10 17 18 12 25 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6118 0 0
2
5.90124e-315 0
0
7 74LS251
144 1023 801 0 14 29
0 38 39 40 41 42 43 44 13 27
28 29 26 45 4
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
45435.4 1
0
7 74LS251
144 1027 699 0 14 29
0 46 47 48 49 50 51 52 14 27
28 29 26 53 5
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6357 0 0
2
45435.4 2
0
7 74LS251
144 1027 599 0 14 29
0 54 55 56 57 58 59 60 15 27
28 29 26 61 6
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
319 0 0
2
45435.4 3
0
7 74LS251
144 1027 492 0 14 29
0 62 63 64 65 66 67 68 16 27
28 29 26 69 7
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3976 0 0
2
45435.4 4
0
7 74LS251
144 1028 389 0 14 29
0 70 71 72 73 74 75 76 17 27
28 29 26 77 8
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
45435.4 5
0
7 74LS251
144 1034 287 0 14 29
0 78 79 80 81 82 83 84 18 27
28 29 26 85 9
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
523 0 0
2
45435.4 6
0
7 74LS251
144 1033 187 0 14 29
0 86 87 88 89 90 91 92 12 27
28 29 26 93 10
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6748 0 0
2
45435.4 7
0
8 Hex Key~
166 1115 33 0 11 12
0 29 28 27 94 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
6901 0 0
2
45435.4 8
0
7 74LS251
144 1033 94 0 14 29
0 95 96 97 98 99 100 101 25 27
28 29 26 102 11
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
842 0 0
2
45435.4 9
0
12 Hex Display~
7 1859 45 0 18 19
10 4 5 6 7 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3277 0 0
2
45435.4 10
0
8 Hex Key~
166 15 40 0 11 12
0 23 24 30 25 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4212 0 0
2
45435.4 11
0
6 74136~
219 89 163 0 3 22
0 30 25 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4720 0 0
2
45435.4 12
0
12 Hex Display~
7 1799 42 0 18 19
10 8 9 10 11 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5551 0 0
2
45435.4 13
0
6 74136~
219 138 193 0 3 22
0 12 24 18
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6986 0 0
2
45435.4 14
0
8 Hex Key~
166 52 42 0 11 12
0 19 20 21 22 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8745 0 0
2
45435.4 15
0
80
1 6 3 0 0 8320 0 1 4 0 0 3
439 589
491 589
491 527
1 9 2 0 0 4240 0 3 4 0 0 2
482 388
482 449
14 1 4 0 0 8192 0 20 5 0 0 3
1055 837
1417 837
1417 52
14 1 5 0 0 8192 0 21 6 0 0 3
1059 735
1382 735
1382 42
14 1 6 0 0 8192 0 22 7 0 0 3
1059 635
1354 635
1354 41
14 1 7 0 0 8192 0 23 8 0 0 3
1059 528
1332 528
1332 41
14 1 8 0 0 8192 0 24 9 0 0 3
1060 425
1298 425
1298 45
14 1 9 0 0 8192 0 25 10 0 0 3
1066 323
1273 323
1273 49
14 1 10 0 0 4096 0 26 11 0 0 3
1065 223
1250 223
1250 51
14 1 11 0 0 4096 0 28 12 0 0 3
1065 130
1215 130
1215 52
14 1 4 0 0 4224 0 20 29 0 0 3
1055 837
1868 837
1868 69
14 2 5 0 0 4224 0 21 29 0 0 3
1059 735
1862 735
1862 69
14 3 6 0 0 4224 0 22 29 0 0 3
1059 635
1856 635
1856 69
14 4 7 0 0 4224 0 23 29 0 0 3
1059 528
1850 528
1850 69
8 3 12 0 0 12416 0 26 31 0 0 4
1001 223
631 223
631 163
122 163
3 8 13 0 0 8320 0 13 20 0 0 4
418 355
607 355
607 837
991 837
8 3 14 0 0 8320 0 21 14 0 0 4
995 735
600 735
600 331
368 331
3 8 15 0 0 12416 0 15 22 0 0 4
317 295
594 295
594 635
995 635
3 8 16 0 0 12416 0 16 23 0 0 4
270 266
588 266
588 528
995 528
8 3 17 0 0 12416 0 24 17 0 0 4
996 425
617 425
617 225
219 225
3 8 18 0 0 4224 0 33 25 0 0 4
171 193
624 193
624 323
1002 323
3 1 13 0 0 0 0 13 18 0 0 3
418 355
594 355
594 51
2 1 19 0 0 4224 0 13 34 0 0 3
369 364
61 364
61 66
3 1 14 0 0 0 0 14 13 0 0 4
368 331
366 331
366 346
369 346
3 2 14 0 0 0 0 14 18 0 0 3
368 331
588 331
588 51
2 2 20 0 0 8320 0 14 34 0 0 3
319 340
55 340
55 66
3 1 15 0 0 0 0 15 14 0 0 3
317 295
317 322
319 322
3 3 15 0 0 0 0 15 18 0 0 3
317 295
582 295
582 51
2 3 21 0 0 8320 0 15 34 0 0 3
268 304
49 304
49 66
3 1 16 0 0 0 0 16 15 0 0 3
270 266
268 266
268 286
3 4 16 0 0 0 0 16 18 0 0 3
270 266
576 266
576 51
4 2 22 0 0 4224 0 34 16 0 0 3
43 66
43 275
221 275
3 1 17 0 0 0 0 17 16 0 0 4
219 225
220 225
220 257
221 257
3 1 17 0 0 0 0 17 19 0 0 3
219 225
542 225
542 52
1 2 23 0 0 4224 0 30 17 0 0 3
24 64
24 234
170 234
3 1 18 0 0 0 0 33 17 0 0 4
171 193
169 193
169 216
170 216
3 2 18 0 0 0 0 33 19 0 0 3
171 193
536 193
536 52
2 2 24 0 0 4224 0 30 33 0 0 3
18 64
18 202
122 202
3 3 12 0 0 0 0 31 19 0 0 3
122 163
530 163
530 52
4 4 25 0 0 8192 0 30 19 0 0 4
6 64
6 130
524 130
524 52
12 1 26 0 0 8320 0 20 2 0 0 3
1061 801
1160 801
1160 34
12 1 26 0 0 0 0 21 2 0 0 3
1065 699
1160 699
1160 34
12 1 26 0 0 0 0 22 2 0 0 3
1065 599
1160 599
1160 34
12 1 26 0 0 0 0 23 2 0 0 3
1065 492
1160 492
1160 34
12 1 26 0 0 0 0 24 2 0 0 3
1066 389
1160 389
1160 34
12 1 26 0 0 0 0 25 2 0 0 3
1072 287
1160 287
1160 34
12 1 26 0 0 0 0 26 2 0 0 3
1071 187
1160 187
1160 34
1 12 26 0 0 0 0 2 28 0 0 3
1160 34
1160 94
1071 94
14 1 8 0 0 4224 0 24 32 0 0 3
1060 425
1808 425
1808 66
14 2 9 0 0 4224 0 25 32 0 0 3
1066 323
1802 323
1802 66
14 3 10 0 0 4224 0 26 32 0 0 3
1065 223
1796 223
1796 66
14 4 11 0 0 4224 0 28 32 0 0 3
1065 130
1790 130
1790 66
9 3 27 0 0 8192 0 22 27 0 0 3
1059 572
1112 572
1112 57
9 3 27 0 0 8192 0 21 27 0 0 3
1059 672
1112 672
1112 57
3 9 27 0 0 4224 0 27 20 0 0 3
1112 57
1112 774
1055 774
10 2 28 0 0 8320 0 20 27 0 0 3
1055 783
1118 783
1118 57
10 2 28 0 0 0 0 21 27 0 0 3
1059 681
1118 681
1118 57
2 10 28 0 0 0 0 27 22 0 0 3
1118 57
1118 581
1059 581
11 1 29 0 0 8320 0 20 27 0 0 3
1055 792
1124 792
1124 57
11 1 29 0 0 0 0 21 27 0 0 3
1059 690
1124 690
1124 57
11 1 29 0 0 0 0 22 27 0 0 3
1059 590
1124 590
1124 57
9 3 27 0 0 0 0 23 27 0 0 3
1059 465
1112 465
1112 57
9 3 27 0 0 0 0 24 27 0 0 3
1060 362
1112 362
1112 57
2 10 28 0 0 0 0 27 23 0 0 3
1118 57
1118 474
1059 474
2 10 28 0 0 0 0 27 24 0 0 3
1118 57
1118 371
1060 371
11 1 29 0 0 0 0 23 27 0 0 3
1059 483
1124 483
1124 57
1 11 29 0 0 0 0 27 24 0 0 3
1124 57
1124 380
1060 380
4 8 25 0 0 8320 0 30 28 0 0 3
6 64
6 130
1001 130
1 11 29 0 0 0 0 27 25 0 0 3
1124 57
1124 278
1066 278
10 2 28 0 0 0 0 25 27 0 0 3
1066 269
1118 269
1118 57
3 9 27 0 0 0 0 27 25 0 0 3
1112 57
1112 260
1066 260
11 1 29 0 0 0 0 26 27 0 0 3
1065 178
1124 178
1124 57
2 10 28 0 0 0 0 27 26 0 0 3
1118 57
1118 169
1065 169
9 3 27 0 0 0 0 26 27 0 0 3
1065 160
1112 160
1112 57
3 9 27 0 0 0 0 27 28 0 0 3
1112 57
1112 67
1065 67
2 10 28 0 0 0 0 27 28 0 0 3
1118 57
1118 76
1065 76
1 11 29 0 0 0 0 27 28 0 0 3
1124 57
1124 85
1065 85
3 1 30 0 0 4224 0 30 31 0 0 3
12 64
12 154
73 154
4 2 25 0 0 0 0 30 31 0 0 3
6 64
6 172
73 172
3 1 12 0 0 0 0 31 33 0 0 2
122 163
122 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
