CircuitMaker Text
5.6
Probes: 1
KPD1_3
Transient Analysis
0 203 83 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
950 130 30 200 10
244 80 1598 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
921 80 1598 839
42991634 0
0
6 Title:
5 Name:
0
0
0
37
7 Ground~
168 1488 466 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6652 0 0
2
5.90125e-315 0
0
6 74LS48
188 295 623 0 14 29
0 36 37 38 39 40 41 42 43 44
45 46 47 48 49
0
0 0 4832 0
6 74LS48
-21 -60 21 -52
3 U14
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4281 0 0
2
5.90125e-315 0
0
6 74LS48
188 295 502 0 14 29
0 50 51 52 53 54 55 56 57 58
59 60 61 62 63
0
0 0 4832 0
6 74LS48
-21 -60 21 -52
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6847 0 0
2
5.90125e-315 5.26354e-315
0
7 74LS151
20 929 915 0 14 29
0 64 65 66 67 68 28 2 29 2
2 13 12 4 69
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
3 U12
55 -5 76 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
6543 0 0
2
5.90125e-315 5.30499e-315
0
7 74LS151
20 929 1013 0 14 29
0 70 71 72 73 74 21 2 21 2
2 13 12 14 75
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
3 U11
55 -5 76 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7168 0 0
2
5.90125e-315 5.32571e-315
0
7 74LS151
20 931 719 0 14 29
0 76 77 78 79 80 26 2 31 2
2 13 12 8 81
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
3 U10
55 -5 76 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3828 0 0
2
5.90125e-315 5.34643e-315
0
7 74LS151
20 929 814 0 14 29
0 82 83 84 85 86 27 2 30 2
2 13 12 9 87
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
2 U9
56 -5 70 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
955 0 0
2
5.90125e-315 5.3568e-315
0
7 74LS151
20 933 526 0 14 29
0 88 89 90 91 92 24 2 33 2
2 13 12 6 93
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
2 U8
56 -5 70 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7782 0 0
2
5.90125e-315 5.36716e-315
0
7 74LS151
20 932 624 0 14 29
0 94 95 96 97 98 25 2 32 2
2 13 12 7 99
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
2 U7
56 -5 70 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
824 0 0
2
5.90125e-315 5.37752e-315
0
7 74LS151
20 933 433 0 14 29
0 100 101 102 103 104 23 2 34 2
2 13 12 5 105
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
2 U6
56 -5 70 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
6983 0 0
2
5.90125e-315 5.38788e-315
0
7 74LS151
20 935 342 0 14 29
0 106 107 108 109 110 22 2 35 2
2 13 12 3 111
0
0 0 4832 90
7 74LS151
-24 -60 25 -52
2 U5
56 -5 70 3
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3185 0 0
2
5.90125e-315 5.39306e-315
0
9 CA 7-Seg~
184 1381 116 0 18 19
10 3 2 2 3 3 3 10 10 112
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
-19 -58 16 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4213 0 0
2
5.90125e-315 5.39824e-315
0
9 CA 7-Seg~
184 1325 116 0 18 19
10 5 2 2 5 5 5 10 10 113
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9765 0 0
2
5.90125e-315 5.40342e-315
0
9 CA 7-Seg~
184 1269 116 0 18 19
10 6 2 2 6 6 6 10 10 114
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8986 0 0
2
5.90125e-315 5.4086e-315
0
9 CA 7-Seg~
184 1213 116 0 18 19
10 7 2 2 7 7 7 10 10 115
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3273 0 0
2
5.90125e-315 5.41378e-315
0
9 CA 7-Seg~
184 1157 116 0 18 19
10 8 2 2 8 8 8 10 10 116
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5636 0 0
2
5.90125e-315 5.41896e-315
0
9 CA 7-Seg~
184 1101 116 0 18 19
10 9 2 2 9 9 9 10 10 117
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP6
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
327 0 0
2
5.90125e-315 5.42414e-315
0
9 CA 7-Seg~
184 1044 116 0 18 19
10 4 2 2 4 4 4 10 10 118
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP8
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9233 0 0
2
5.90125e-315 5.42933e-315
0
9 CA 7-Seg~
184 988 116 0 18 19
10 14 2 2 14 14 14 10 10 119
0 0 0 0 0 0 1 1 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP7
-16 -58 19 -50
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3875 0 0
2
5.90125e-315 5.43192e-315
0
9 2-In XOR~
219 718 181 0 3 22
0 15 11 35
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U1A
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
9991 0 0
2
5.90125e-315 5.43451e-315
0
9 2-In XOR~
219 718 280 0 3 22
0 17 18 32
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U1C
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3221 0 0
2
5.90125e-315 5.4371e-315
0
9 2-In XOR~
219 718 247 0 3 22
0 16 17 33
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U1D
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8874 0 0
2
5.90125e-315 5.43969e-315
0
9 2-In XOR~
219 718 214 0 3 22
0 11 16 34
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U1B
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7400 0 0
2
5.90125e-315 5.44228e-315
0
9 2-In XOR~
219 718 313 0 3 22
0 18 20 31
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U2A
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3623 0 0
2
5.90125e-315 5.44487e-315
0
9 2-In XOR~
219 718 346 0 3 22
0 20 19 30
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U2B
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3311 0 0
2
5.90125e-315 5.44746e-315
0
9 2-In XOR~
219 718 379 0 3 22
0 19 21 29
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U2C
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5736 0 0
2
5.90125e-315 5.45005e-315
0
2 +V
167 1487 60 0 1 3
0 10
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3143 0 0
2
5.90125e-315 5.45264e-315
0
9 2-In XOR~
219 723 957 0 3 22
0 18 27 26
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3C
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5835 0 0
2
5.90125e-315 5.45782e-315
0
9 2-In XOR~
219 723 825 0 3 22
0 15 23 22
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U4C
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
5108 0 0
2
5.90125e-315 5.46041e-315
0
9 2-In XOR~
219 723 924 0 3 22
0 17 26 25
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U4B
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3320 0 0
2
5.90125e-315 5.463e-315
0
9 2-In XOR~
219 723 891 0 3 22
0 16 25 24
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U4A
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
523 0 0
2
5.90125e-315 5.46559e-315
0
9 2-In XOR~
219 723 858 0 3 22
0 11 24 23
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3D
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3557 0 0
2
5.90125e-315 5.46818e-315
0
9 2-In XOR~
219 723 990 0 3 22
0 20 28 27
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3B
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7246 0 0
2
5.90125e-315 5.47077e-315
0
9 2-In XOR~
219 723 1023 0 3 22
0 19 21 28
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3A
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3916 0 0
2
5.90125e-315 5.47207e-315
0
8 Hex Key~
166 47 49 0 11 12
0 12 13 120 121 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
614 0 0
2
45437.8 0
0
8 Hex Key~
166 85 49 0 11 12
0 18 20 19 21 0 0 0 0 0
15 70
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8494 0 0
2
45437.8 1
0
8 Hex Key~
166 126 49 0 11 12
0 15 11 16 17 0 0 0 0 0
15 70
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
774 0 0
2
45437.8 2
0
156
4 0 0 0 0 0 0 2 0 0 72 2
263 614
94 614
3 0 0 0 0 0 0 2 0 0 74 2
263 605
88 605
2 0 0 0 0 0 0 2 0 0 73 2
263 596
82 596
1 0 0 0 0 0 0 2 0 0 97 2
263 587
76 587
4 0 0 0 0 0 0 3 0 0 69 2
263 493
135 493
3 0 0 0 0 0 0 3 0 0 36 2
263 484
129 484
2 0 0 0 0 0 0 3 0 0 70 2
263 475
123 475
1 0 0 0 0 0 0 3 0 0 71 2
263 466
118 466
5 0 3 0 0 4096 0 12 0 0 21 2
1384 152
1384 167
0 4 3 0 0 0 0 0 12 21 0 2
1378 167
1378 152
0 1 3 0 0 0 0 0 12 21 0 2
1360 167
1360 152
0 7 2 0 0 8192 0 0 11 52 0 3
1000 376
1000 374
968 374
7 0 2 0 0 8192 0 10 0 0 52 3
966 465
966 468
1000 468
7 0 2 0 0 0 0 8 0 0 52 3
966 558
966 563
1000 563
7 0 2 0 0 8192 0 9 0 0 52 3
965 656
965 659
1000 659
7 0 2 0 0 8192 0 6 0 0 52 3
964 751
964 755
1000 755
7 0 2 0 0 8192 0 7 0 0 52 3
962 846
962 850
1000 850
0 7 2 0 0 0 0 0 4 52 0 3
1000 952
962 952
962 947
0 7 2 0 0 4096 0 0 5 52 0 4
1000 961
1000 1051
962 1051
962 1045
0 13 4 0 0 12416 0 0 4 129 0 6
1023 165
1023 286
1007 286
1007 865
962 865
962 883
6 13 3 0 0 16528 0 12 11 0 0 8
1390 152
1390 167
1360 167
1360 262
1019 262
1019 298
968 298
968 310
0 13 5 0 0 8320 0 0 10 117 0 6
1304 167
1304 266
1017 266
1017 390
966 390
966 401
0 9 2 0 0 0 0 0 5 52 0 3
918 961
908 961
908 975
0 9 2 0 0 0 0 0 4 51 0 3
917 859
908 859
908 877
0 9 2 0 0 0 0 0 7 50 0 3
917 763
908 763
908 776
0 9 2 0 0 0 0 0 6 49 0 3
919 667
910 667
910 681
0 9 2 0 0 0 0 0 9 48 0 3
920 572
911 572
911 586
0 9 2 0 0 0 0 0 8 47 0 3
921 476
912 476
912 488
0 9 2 0 0 0 0 0 10 46 0 3
921 384
912 384
912 395
0 9 2 0 0 0 0 0 11 44 0 3
923 292
914 292
914 304
0 13 6 0 0 8320 0 0 8 120 0 6
1248 166
1248 270
1015 270
1015 482
966 482
966 494
0 13 7 0 0 12416 0 0 9 123 0 6
1192 165
1192 274
1013 274
1013 578
965 578
965 592
0 13 8 0 0 12416 0 0 6 126 0 6
1136 168
1136 278
1011 278
1011 673
964 673
964 687
0 13 9 0 0 12416 0 0 7 114 0 6
1080 164
1080 282
1009 282
1009 769
962 769
962 782
8 0 10 0 0 4096 0 17 0 0 156 2
1122 152
1122 254
1 0 11 0 0 8320 0 32 0 0 77 3
707 849
129 849
129 205
8 0 10 0 0 0 0 12 0 0 156 2
1402 152
1402 254
8 0 10 0 0 0 0 13 0 0 156 2
1346 152
1346 254
8 0 10 0 0 0 0 14 0 0 156 2
1290 152
1290 254
8 0 10 0 0 0 0 15 0 0 156 2
1234 152
1234 254
8 0 10 0 0 0 0 16 0 0 156 2
1178 152
1178 254
8 0 10 0 0 0 0 18 0 0 156 2
1065 152
1065 254
8 0 10 0 0 0 0 19 0 0 156 2
1009 152
1009 254
10 0 2 0 0 0 0 11 0 0 52 3
923 310
923 292
1000 292
12 0 12 0 0 8192 0 10 0 0 67 3
939 401
939 388
992 388
10 0 2 0 0 0 0 10 0 0 52 3
921 401
921 384
1000 384
10 0 2 0 0 0 0 8 0 0 52 3
921 494
921 476
1000 476
10 0 2 0 0 0 0 9 0 0 52 3
920 592
920 572
1000 572
10 0 2 0 0 0 0 6 0 0 52 3
919 687
919 667
1000 667
10 0 2 0 0 0 0 7 0 0 52 3
917 782
917 763
1000 763
10 0 2 0 0 0 0 4 0 0 52 3
917 883
917 859
1000 859
0 10 2 0 0 4224 0 0 5 148 0 4
1000 258
1000 961
917 961
917 981
11 0 13 0 0 8192 0 5 0 0 66 3
926 981
926 963
994 963
12 0 12 0 0 8192 0 5 0 0 67 3
935 981
935 965
992 965
11 0 13 0 0 0 0 4 0 0 66 3
926 883
926 861
994 861
12 0 12 0 0 0 0 4 0 0 67 3
935 883
935 863
992 863
11 0 13 0 0 0 0 7 0 0 66 3
926 782
926 765
994 765
12 0 12 0 0 0 0 7 0 0 67 3
935 782
935 767
992 767
11 0 13 0 0 0 0 6 0 0 66 3
928 687
928 669
994 669
11 0 13 0 0 0 0 9 0 0 66 3
929 592
929 574
994 574
11 0 13 0 0 0 0 8 0 0 66 3
930 494
930 478
994 478
12 0 12 0 0 0 0 6 0 0 67 3
937 687
937 671
992 671
12 0 12 0 0 0 0 9 0 0 67 3
938 592
938 576
992 576
12 0 12 0 0 0 0 8 0 0 67 3
939 494
939 480
992 480
0 11 13 0 0 0 0 0 10 66 0 3
994 386
930 386
930 401
2 11 13 0 0 4224 0 35 11 0 0 6
50 73
50 1081
994 1081
994 294
932 294
932 310
1 12 12 0 0 4224 0 35 11 0 0 6
56 73
56 1075
992 1075
992 296
941 296
941 310
0 13 14 0 0 12416 0 0 5 132 0 6
967 165
967 290
1005 290
1005 967
962 967
962 981
0 1 15 0 0 4224 0 0 29 75 0 3
135 172
135 816
707 816
0 1 16 0 0 4224 0 0 31 79 0 3
123 238
123 882
707 882
0 1 17 0 0 4224 0 0 30 81 0 3
118 271
118 915
707 915
0 1 18 0 0 4224 0 0 28 83 0 3
94 304
94 948
707 948
0 1 19 0 0 4224 0 0 34 87 0 3
82 370
82 1014
707 1014
0 1 20 0 0 4224 0 0 33 85 0 3
88 337
88 981
707 981
1 1 15 0 0 0 0 20 37 0 0 3
702 172
135 172
135 73
2 0 11 0 0 0 0 20 0 0 77 2
702 190
129 190
1 2 11 0 0 0 0 23 37 0 0 3
702 205
129 205
129 73
2 0 16 0 0 0 0 23 0 0 79 2
702 223
123 223
1 3 16 0 0 0 0 22 37 0 0 3
702 238
123 238
123 73
2 0 17 0 0 0 0 22 0 0 81 2
702 256
117 256
1 4 17 0 0 0 0 21 37 0 0 3
702 271
117 271
117 73
2 0 18 0 0 0 0 21 0 0 83 2
702 289
94 289
1 1 18 0 0 0 0 24 36 0 0 3
702 304
94 304
94 73
2 0 20 0 0 0 0 24 0 0 85 2
702 322
88 322
1 2 20 0 0 0 0 25 36 0 0 3
702 337
88 337
88 73
2 0 19 0 0 0 0 25 0 0 87 2
702 355
82 355
1 3 19 0 0 0 0 26 36 0 0 3
702 370
82 370
82 73
2 0 21 0 0 4096 0 26 0 0 98 2
702 388
76 388
2 0 21 0 0 4096 0 34 0 0 97 2
707 1032
76 1032
6 3 22 0 0 12416 0 11 29 0 0 5
959 374
959 382
857 382
857 825
756 825
6 3 23 0 0 12416 0 10 32 0 0 5
957 465
957 474
859 474
859 858
756 858
6 3 24 0 0 12416 0 8 31 0 0 5
957 558
957 570
861 570
861 891
756 891
6 3 25 0 0 12416 0 9 30 0 0 5
956 656
956 665
863 665
863 924
756 924
6 3 26 0 0 12416 0 6 28 0 0 5
955 751
955 761
865 761
865 957
756 957
6 3 27 0 0 12416 0 7 33 0 0 5
953 846
953 857
867 857
867 990
756 990
6 3 28 0 0 16512 0 4 34 0 0 5
953 947
953 959
869 959
869 1023
756 1023
0 6 21 0 0 8320 0 0 5 98 0 4
76 409
76 1057
953 1057
953 1045
4 8 21 0 0 0 0 36 5 0 0 6
76 73
76 409
874 409
874 1055
971 1055
971 1045
8 3 29 0 0 12416 0 4 26 0 0 5
971 947
971 957
876 957
876 379
751 379
8 3 30 0 0 12416 0 7 25 0 0 5
971 846
971 855
878 855
878 346
751 346
8 3 31 0 0 12416 0 6 24 0 0 5
973 751
973 759
880 759
880 313
751 313
8 3 32 0 0 12416 0 9 21 0 0 5
974 656
974 663
882 663
882 280
751 280
8 3 33 0 0 12416 0 8 22 0 0 5
975 558
975 568
884 568
884 247
751 247
8 3 34 0 0 12416 0 10 23 0 0 5
975 465
975 472
886 472
886 214
751 214
8 3 35 0 0 12416 0 11 20 0 0 5
977 374
977 380
888 380
888 181
751 181
3 2 23 0 0 0 0 32 29 0 0 5
756 858
756 841
677 841
677 834
707 834
3 2 24 0 0 0 0 31 32 0 0 5
756 891
756 874
675 874
675 867
707 867
3 2 25 0 0 0 0 30 31 0 0 5
756 924
756 906
675 906
675 900
707 900
3 2 26 0 0 0 0 28 30 0 0 5
756 957
756 940
677 940
677 933
707 933
3 2 27 0 0 0 0 33 28 0 0 5
756 990
756 973
676 973
676 966
707 966
3 2 28 0 0 0 0 34 33 0 0 5
756 1023
756 1006
675 1006
675 999
707 999
0 6 9 0 0 0 0 0 17 113 0 3
1104 158
1110 158
1110 152
0 5 9 0 0 0 0 0 17 114 0 3
1098 164
1104 164
1104 152
1 4 9 0 0 0 0 17 17 0 0 4
1080 152
1080 164
1098 164
1098 152
0 6 5 0 0 0 0 0 13 116 0 3
1328 167
1334 167
1334 152
0 5 5 0 0 0 0 0 13 117 0 3
1321 167
1328 167
1328 152
1 4 5 0 0 0 0 13 13 0 0 4
1304 152
1304 167
1322 167
1322 152
0 6 6 0 0 0 0 0 14 119 0 3
1272 166
1278 166
1278 152
0 5 6 0 0 0 0 0 14 120 0 3
1266 166
1272 166
1272 152
1 4 6 0 0 0 0 14 14 0 0 4
1248 152
1248 166
1266 166
1266 152
0 6 7 0 0 0 0 0 15 122 0 3
1216 165
1222 165
1222 152
0 5 7 0 0 0 0 0 15 123 0 3
1210 165
1216 165
1216 152
1 4 7 0 0 0 0 15 15 0 0 4
1192 152
1192 165
1210 165
1210 152
0 6 8 0 0 0 0 0 16 125 0 3
1160 168
1166 168
1166 152
0 5 8 0 0 0 0 0 16 126 0 3
1154 168
1160 168
1160 152
1 4 8 0 0 0 0 16 16 0 0 4
1136 152
1136 168
1154 168
1154 152
0 6 4 0 0 0 0 0 18 128 0 3
1047 165
1053 165
1053 152
0 5 4 0 0 0 0 0 18 129 0 3
1040 165
1047 165
1047 152
1 4 4 0 0 0 0 18 18 0 0 4
1023 152
1023 165
1041 165
1041 152
0 6 14 0 0 0 0 0 19 131 0 3
991 159
997 159
997 152
0 5 14 0 0 0 0 0 19 132 0 3
985 165
991 165
991 152
1 4 14 0 0 0 0 19 19 0 0 4
967 152
967 165
985 165
985 152
3 0 2 0 0 0 0 12 0 0 148 2
1372 152
1372 258
2 0 2 0 0 0 0 12 0 0 148 2
1366 152
1366 258
3 0 2 0 0 0 0 13 0 0 148 2
1316 152
1316 258
2 0 2 0 0 0 0 13 0 0 148 2
1310 152
1310 258
3 0 2 0 0 0 0 14 0 0 148 2
1260 152
1260 258
2 0 2 0 0 0 0 14 0 0 148 2
1254 152
1254 258
3 0 2 0 0 0 0 15 0 0 148 2
1204 152
1204 258
2 0 2 0 0 0 0 15 0 0 148 2
1198 152
1198 258
3 0 2 0 0 0 0 16 0 0 148 2
1148 152
1148 258
2 0 2 0 0 0 0 16 0 0 148 2
1142 152
1142 258
3 0 2 0 0 0 0 17 0 0 148 2
1092 152
1092 258
2 0 2 0 0 0 0 17 0 0 148 2
1086 152
1086 258
3 0 2 0 0 0 0 18 0 0 148 2
1035 152
1035 258
2 0 2 0 0 0 0 18 0 0 148 2
1029 152
1029 258
3 0 2 0 0 0 0 19 0 0 148 2
979 152
979 258
1 2 2 0 0 0 0 1 19 0 0 4
1488 460
1488 258
973 258
973 152
7 0 10 0 0 0 0 12 0 0 156 2
1396 152
1396 254
7 0 10 0 0 0 0 13 0 0 156 2
1340 152
1340 254
7 0 10 0 0 0 0 14 0 0 156 2
1284 152
1284 254
7 0 10 0 0 0 0 15 0 0 156 2
1228 152
1228 254
7 0 10 0 0 0 0 16 0 0 156 2
1172 152
1172 254
7 0 10 0 0 0 0 17 0 0 156 2
1116 152
1116 254
7 0 10 0 0 0 0 18 0 0 156 2
1059 152
1059 254
1 7 10 0 0 8320 0 27 19 0 0 4
1487 69
1487 254
1003 254
1003 152
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
