CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
34
14 Logic Display~
6 1153 24 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
45435.5 0
0
14 Logic Display~
6 1121 27 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
45435.5 0
0
14 Logic Display~
6 1091 27 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
45435.5 0
0
14 Logic Display~
6 1061 25 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
45435.5 0
0
14 Logic Display~
6 1031 27 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
45435.5 0
0
14 Logic Display~
6 999 27 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
45435.5 0
0
14 Logic Display~
6 969 29 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
45435.5 0
0
14 Logic Display~
6 941 31 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 1 0 0
1 L
34 0 0
2
45435.5 0
0
6 74136~
219 140 715 0 3 22
0 18 17 2
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
969 0 0
2
45435.5 0
0
6 74136~
219 134 671 0 3 22
0 19 18 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8402 0 0
2
45435.5 0
0
6 74136~
219 137 623 0 3 22
0 20 19 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3751 0 0
2
45435.5 0
0
6 74136~
219 138 565 0 3 22
0 21 20 5
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4292 0 0
2
45435.5 0
0
6 74136~
219 140 516 0 3 22
0 22 21 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6118 0 0
2
45435.5 0
0
6 74136~
219 138 469 0 3 22
0 23 23 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
34 0 0
2
45435.5 0
0
6 74136~
219 136 417 0 3 22
0 9 23 8
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
6357 0 0
2
45435.5 0
0
7 Ground~
168 1450 261 0 1 3
0 24
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
319 0 0
2
5.90124e-315 0
0
9 CC 7-Seg~
183 1558 431 0 18 19
10 25 26 27 28 29 30 31 32 33
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3976 0 0
2
5.90124e-315 0
0
14 Logic Display~
6 811 37 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
45435.5 0
0
14 Logic Display~
6 773 35 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
45435.5 1
0
14 Logic Display~
6 742 36 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
45435.5 2
0
14 Logic Display~
6 705 38 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
45435.5 3
0
14 Logic Display~
6 670 39 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
45435.5 4
0
14 Logic Display~
6 636 39 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
45435.5 5
0
14 Logic Display~
6 601 39 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
45435.5 6
0
14 Logic Display~
6 568 40 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
45435.5 7
0
6 74136~
219 385 355 0 3 22
0 11 17 10
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5551 0 0
2
45435.5 8
0
6 74136~
219 335 326 0 3 22
0 12 18 11
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6986 0 0
2
45435.5 9
0
6 74136~
219 284 295 0 3 22
0 13 19 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8745 0 0
2
45435.5 10
0
6 74136~
219 237 266 0 3 22
0 14 20 13
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9592 0 0
2
45435.5 11
0
6 74136~
219 186 225 0 3 22
0 15 21 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8748 0 0
2
45435.5 12
0
8 Hex Key~
166 15 40 0 11 12
0 21 22 23 9 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7168 0 0
2
5.90124e-315 5.40342e-315
0
6 74136~
219 89 163 0 3 22
0 23 9 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
631 0 0
2
5.90124e-315 5.4086e-315
0
6 74136~
219 138 193 0 3 22
0 16 22 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9466 0 0
2
5.90124e-315 5.41896e-315
0
8 Hex Key~
166 52 42 0 11 12
0 17 18 19 20 0 0 0 0 0
15 70
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3266 0 0
2
5.90124e-315 5.42414e-315
0
44
1 3 2 0 0 8320 0 1 9 0 0 3
1153 42
1153 715
173 715
3 1 3 0 0 4224 0 10 2 0 0 3
167 671
1121 671
1121 45
3 1 4 0 0 4224 0 11 3 0 0 3
170 623
1091 623
1091 45
3 1 5 0 0 4224 0 12 4 0 0 3
171 565
1061 565
1061 43
3 1 6 0 0 4224 0 13 5 0 0 3
173 516
1031 516
1031 45
3 1 7 0 0 4224 0 14 6 0 0 3
171 469
999 469
999 45
3 1 8 0 0 4224 0 15 7 0 0 3
169 417
969 417
969 47
4 1 9 0 0 8336 0 31 8 0 0 4
6 64
6 387
941 387
941 49
3 1 10 0 0 4224 0 26 18 0 0 3
418 355
811 355
811 55
3 1 11 0 0 4224 0 27 19 0 0 3
368 326
773 326
773 53
3 1 12 0 0 4224 0 28 20 0 0 3
317 295
742 295
742 54
3 1 13 0 0 4224 0 29 21 0 0 3
270 266
705 266
705 56
3 1 14 0 0 4224 0 30 22 0 0 3
219 225
670 225
670 57
3 1 15 0 0 4224 0 33 23 0 0 3
171 193
636 193
636 57
3 1 16 0 0 4224 0 32 24 0 0 3
122 163
601 163
601 57
4 1 9 0 0 0 0 31 25 0 0 4
6 64
6 71
568 71
568 58
1 2 17 0 0 4224 0 34 9 0 0 3
61 66
61 724
124 724
2 1 18 0 0 4224 0 34 9 0 0 3
55 66
55 706
124 706
2 2 18 0 0 0 0 34 10 0 0 3
55 66
55 680
118 680
3 1 19 0 0 4224 0 34 10 0 0 3
49 66
49 662
118 662
3 2 19 0 0 0 0 34 11 0 0 3
49 66
49 632
121 632
4 1 20 0 0 4224 0 34 11 0 0 3
43 66
43 614
121 614
4 2 20 0 0 0 0 34 12 0 0 3
43 66
43 574
122 574
1 1 21 0 0 8320 0 12 31 0 0 3
122 556
24 556
24 64
1 2 21 0 0 0 0 31 13 0 0 3
24 64
24 525
124 525
2 1 22 0 0 4224 0 31 13 0 0 3
18 64
18 507
124 507
3 2 23 0 0 4224 0 31 14 0 0 3
12 64
12 478
122 478
3 1 23 0 0 0 0 31 14 0 0 3
12 64
12 460
122 460
3 2 23 0 0 0 0 31 15 0 0 3
12 64
12 426
120 426
4 1 9 0 0 0 0 31 15 0 0 3
6 64
6 408
120 408
2 1 17 0 0 128 0 26 34 0 0 3
369 364
61 364
61 66
3 1 11 0 0 0 0 27 26 0 0 4
368 326
366 326
366 346
369 346
2 2 18 0 0 128 0 27 34 0 0 3
319 335
55 335
55 66
3 1 12 0 0 0 0 28 27 0 0 3
317 295
317 317
319 317
2 3 19 0 0 128 0 28 34 0 0 3
268 304
49 304
49 66
3 1 13 0 0 0 0 29 28 0 0 3
270 266
268 266
268 286
4 2 20 0 0 128 0 34 29 0 0 3
43 66
43 275
221 275
3 1 14 0 0 0 0 30 29 0 0 4
219 225
220 225
220 257
221 257
1 2 21 0 0 128 0 31 30 0 0 3
24 64
24 234
170 234
3 1 15 0 0 0 0 33 30 0 0 4
171 193
169 193
169 216
170 216
2 2 22 0 0 128 0 31 33 0 0 3
18 64
18 202
122 202
3 1 23 0 0 128 0 31 32 0 0 3
12 64
12 154
73 154
4 2 9 0 0 0 0 31 32 0 0 3
6 64
6 172
73 172
3 1 16 0 0 0 0 32 33 0 0 2
122 163
122 184
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
449 15 550 39
460 24 538 40
13 Grey->Binario
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
831 16 932 40
842 25 920 41
13 Binario->Grey
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
152 429 243 453
164 438 230 454
11 Codificador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
223 192 330 216
234 201 318 217
14 DE_Codificador
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
