CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
110
13 Logic Switch~
5 790 2347 0 1 11
0 20
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 1160 22 0 1 11
0 104
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90125e-315 5.26354e-315
0
9 Inverter~
13 183 927 0 2 22
0 6 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 29 0
1 U
3124 0 0
2
45438.7 0
0
9 Inverter~
13 120 1009 0 2 22
0 5 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 29 0
1 U
3421 0 0
2
45438.7 0
0
9 Inverter~
13 163 1000 0 2 22
0 6 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 29 0
1 U
8157 0 0
2
45438.7 0
0
9 Inverter~
13 203 991 0 2 22
0 7 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 29 0
1 U
5572 0 0
2
45438.7 0
0
5 7415~
219 349 1000 0 4 22
0 10 9 8 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 8 0
1 U
8901 0 0
2
45438.7 0
0
5 7415~
219 348 927 0 4 22
0 7 11 5 3
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U27C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 22 0
1 U
7361 0 0
2
45438.7 0
0
9 Inverter~
13 215 2268 0 2 22
0 6 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 27 0
1 U
4747 0 0
2
45438.7 0
0
9 Inverter~
13 206 2215 0 2 22
0 7 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 27 0
1 U
972 0 0
2
45438.7 0
0
9 Inverter~
13 220 2172 0 2 22
0 5 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 27 0
1 U
3472 0 0
2
45438.7 0
0
9 2-In AND~
219 402 2259 0 3 22
0 7 21 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
9998 0 0
2
45438.7 0
0
9 2-In AND~
219 345 2224 0 3 22
0 22 6 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
3536 0 0
2
45438.7 0
0
9 2-In AND~
219 394 2181 0 3 22
0 23 6 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
4597 0 0
2
45438.7 0
0
8 4-In OR~
219 562 2173 0 5 22
0 12 26 25 24 13
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 25 0
1 U
3835 0 0
2
45438.7 0
0
9 Inverter~
13 233 2079 0 2 22
0 6 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 27 0
1 U
3670 0 0
2
45438.7 0
0
9 Inverter~
13 233 2027 0 2 22
0 5 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 27 0
1 U
5616 0 0
2
45438.7 0
0
9 Inverter~
13 201 1973 0 2 22
0 6 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 27 0
1 U
9323 0 0
2
45438.7 0
0
9 Inverter~
13 144 1991 0 2 22
0 5 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28F
-14 -18 14 -10
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 23 0
1 U
317 0 0
2
45438.7 0
0
9 2-In AND~
219 371 2070 0 3 22
0 7 29 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
3108 0 0
2
45438.7 0
0
9 2-In AND~
219 367 2018 0 3 22
0 7 30 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
4299 0 0
2
45438.7 0
0
9 2-In AND~
219 309 1982 0 3 22
0 33 32 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
9672 0 0
2
45438.7 0
0
8 4-In OR~
219 554 1976 0 5 22
0 12 31 28 27 14
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 25 0
1 U
7876 0 0
2
45438.7 0
0
9 Inverter~
13 214 1383 0 2 22
0 12 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 23 0
1 U
6369 0 0
2
45438.7 0
0
9 Inverter~
13 242 1374 0 2 22
0 6 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 23 0
1 U
9172 0 0
2
45438.7 0
0
9 Inverter~
13 273 1365 0 2 22
0 5 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 23 0
1 U
7100 0 0
2
45438.7 0
0
5 7415~
219 381 1374 0 4 22
0 37 36 35 38
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U27B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 22 0
1 U
3820 0 0
2
45438.7 0
0
9 4-In AND~
219 414 1784 0 5 22
0 7 40 5 39 34
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U29A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 24 0
1 U
7678 0 0
2
45438.7 0
0
9 Inverter~
13 194 1798 0 2 22
0 12 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 23 0
1 U
961 0 0
2
45438.7 0
0
9 Inverter~
13 130 1750 0 2 22
0 12 43
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 23 0
1 U
3178 0 0
2
45438.7 0
0
9 Inverter~
13 214 1741 0 2 22
0 7 42
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 21 0
1 U
3409 0 0
2
45438.7 0
0
9 Inverter~
13 284 1732 0 2 22
0 5 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 21 0
1 U
3951 0 0
2
45438.7 0
0
9 Inverter~
13 173 1780 0 2 22
0 6 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 21 0
1 U
8885 0 0
2
45438.7 0
0
9 Inverter~
13 169 1828 0 2 22
0 5 45
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 21 0
1 U
3780 0 0
2
45438.7 0
0
9 Inverter~
13 162 1892 0 2 22
0 5 44
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 21 0
1 U
9265 0 0
2
45438.7 0
0
9 2-In AND~
219 382 1883 0 3 22
0 12 44 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
9442 0 0
2
45438.7 0
0
9 2-In AND~
219 425 1837 0 3 22
0 45 6 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
9424 0 0
2
45438.7 0
0
5 7415~
219 441 1741 0 4 22
0 41 42 43 48
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U27A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 22 0
1 U
9968 0 0
2
45438.7 0
0
8 4-In OR~
219 546 1776 0 5 22
0 48 34 47 46 15
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
9281 0 0
2
45438.7 0
0
9 Inverter~
13 142 1685 0 2 22
0 5 49
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 21 0
1 U
8464 0 0
2
45438.7 0
0
9 Inverter~
13 198 1667 0 2 22
0 12 50
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 20 0
1 U
7168 0 0
2
45438.7 0
0
9 Inverter~
13 167 1622 0 2 22
0 7 51
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 20 0
1 U
3171 0 0
2
45438.7 0
0
9 Inverter~
13 90 1613 0 2 22
0 12 52
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 20 0
1 U
4139 0 0
2
45438.7 0
0
9 Inverter~
13 250 1577 0 2 22
0 6 56
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 20 0
1 U
6435 0 0
2
45438.7 0
0
9 Inverter~
13 171 1568 0 2 22
0 7 57
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 20 0
1 U
5283 0 0
2
45438.7 0
0
9 Inverter~
13 221 1534 0 2 22
0 6 59
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 20 0
1 U
6874 0 0
2
45438.7 0
0
8 Hex Key~
166 54 2358 0 11 12
0 12 7 6 5 0 0 0 0 0
2 50
0
0 0 4656 180
0
4 KPD4
20 -2 48 6
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5305 0 0
2
45438.7 0
0
9 Inverter~
13 182 1506 0 2 22
0 5 61
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 14 0
1 U
34 0 0
2
45438.7 0
0
9 Inverter~
13 231 1497 0 2 22
0 6 62
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 14 0
1 U
969 0 0
2
45438.7 0
0
9 Inverter~
13 278 1488 0 2 22
0 7 63
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 14 0
1 U
8402 0 0
2
45438.7 0
0
5 7415~
219 365 1676 0 4 22
0 50 6 49 53
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 19 0
1 U
3751 0 0
2
45438.7 0
0
5 7415~
219 366 1568 0 4 22
0 12 57 56 55
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 19 0
1 U
4292 0 0
2
45438.7 0
0
5 7415~
219 323 1534 0 4 22
0 7 59 5 58
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 19 0
1 U
6118 0 0
2
45438.7 0
0
5 7415~
219 323 1622 0 4 22
0 52 51 6 54
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 15 0
1 U
34 0 0
2
45438.7 0
0
5 7415~
219 363 1497 0 4 22
0 63 62 61 60
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 15 0
1 U
6357 0 0
2
45438.7 0
0
8 2-In OR~
219 524 1528 0 3 22
0 65 64 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
319 0 0
2
45438.7 0
0
8 2-In OR~
219 433 1646 0 3 22
0 54 53 64
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
3976 0 0
2
45438.7 0
0
8 3-In OR~
219 423 1506 0 4 22
0 60 58 55 65
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U22A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 17 0
1 U
7634 0 0
2
45438.7 0
0
9 2-In AND~
219 335 1418 0 3 22
0 68 67 66
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U21B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
523 0 0
2
45438.7 0
0
5 7415~
219 336 1342 0 4 22
0 6 7 70 69
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 15 0
1 U
6748 0 0
2
45438.7 0
0
5 7415~
219 382 1307 0 4 22
0 72 5 6 71
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U17C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 12 0
1 U
6901 0 0
2
45438.7 0
0
9 Inverter~
13 165 1427 0 2 22
0 6 67
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 14 0
1 U
842 0 0
2
45438.7 0
0
9 Inverter~
13 92 1409 0 2 22
0 7 68
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
3277 0 0
2
45438.7 0
0
9 Inverter~
13 145 1351 0 2 22
0 12 70
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
4212 0 0
2
45438.7 0
0
9 Inverter~
13 168 1298 0 2 22
0 12 72
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
4720 0 0
2
45438.7 0
0
8 4-In OR~
219 523 1320 0 5 22
0 71 69 38 66 17
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
5551 0 0
2
45438.7 0
0
9 Inverter~
13 198 1229 0 2 22
0 6 74
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
6986 0 0
2
45438.7 0
0
9 Inverter~
13 160 1211 0 2 22
0 5 75
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
8745 0 0
2
45438.7 0
0
9 2-In AND~
219 384 1220 0 3 22
0 75 74 73
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
9592 0 0
2
45438.7 0
0
9 2-In AND~
219 311 1194 0 3 22
0 6 5 76
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
8748 0 0
2
45438.7 0
0
9 Inverter~
13 97 1170 0 2 22
0 7 77
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
7168 0 0
2
45438.7 0
0
8 4-In OR~
219 568 1174 0 5 22
0 12 77 76 73 18
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
631 0 0
2
45438.7 0
0
7 Ground~
168 990 922 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9466 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 573 1078 0 5 22
0 12 6 3 4 19
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
3266 0 0
2
5.90125e-315 0
0
9 CC 7-Seg~
183 851 1958 0 15 19
10 19 18 17 16 15 14 13 20 2
1 1 1 1 1 1
0
0 0 21104 270
5 REDCC
16 -41 51 -33
5 DISP3
-21 -39 14 -31
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
7693 0 0
2
5.90125e-315 0
0
6 74136~
219 127 769 0 3 22
0 6 5 79
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3723 0 0
2
5.90125e-315 0
0
6 74136~
219 129 719 0 3 22
0 7 6 80
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3440 0 0
2
5.90125e-315 0
0
6 74136~
219 127 667 0 3 22
0 12 7 81
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6263 0 0
2
5.90125e-315 0
0
6 74136~
219 126 612 0 3 22
0 86 12 85
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4900 0 0
2
5.90125e-315 0
0
6 74136~
219 133 564 0 3 22
0 90 86 87
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
8783 0 0
2
5.90125e-315 0
0
6 74136~
219 126 513 0 3 22
0 91 90 88
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3221 0 0
2
5.90125e-315 0
0
6 74136~
219 200 448 0 3 22
0 78 91 89
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3215 0 0
2
5.90125e-315 0
0
14 Logic Display~
6 1417 34 0 1 2
10 96
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
45438.7 0
0
14 Logic Display~
6 1382 24 0 1 2
10 97
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7121 0 0
2
45438.7 1
0
14 Logic Display~
6 1354 23 0 1 2
10 98
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
45438.7 2
0
14 Logic Display~
6 1332 23 0 1 2
10 99
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
45438.7 3
0
14 Logic Display~
6 1298 27 0 1 2
10 100
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
45438.7 4
0
14 Logic Display~
6 1273 31 0 1 2
10 101
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
45438.7 5
0
14 Logic Display~
6 1250 33 0 1 2
10 102
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
45438.7 6
0
14 Logic Display~
6 1215 34 0 1 2
10 103
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
45438.7 7
0
6 74136~
219 385 355 0 3 22
0 83 5 82
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8396 0 0
2
45438.7 8
0
6 74136~
219 335 331 0 3 22
0 84 6 83
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3685 0 0
2
45438.7 9
0
6 74136~
219 284 295 0 3 22
0 92 7 84
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7849 0 0
2
45438.7 10
0
6 74136~
219 237 266 0 3 22
0 93 12 92
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6343 0 0
2
45438.7 11
0
6 74136~
219 186 225 0 3 22
0 94 86 93
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7376 0 0
2
45438.7 12
0
7 74LS251
144 1023 801 0 14 29
0 108 109 110 111 112 82 113 79 105
106 107 104 114 96
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9156 0 0
2
5.90125e-315 5.34643e-315
0
7 74LS251
144 1027 699 0 14 29
0 115 116 117 118 119 83 120 80 105
106 107 104 121 97
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5776 0 0
2
5.90125e-315 5.3568e-315
0
7 74LS251
144 1027 599 0 14 29
0 122 123 124 125 126 84 127 81 105
106 107 104 128 98
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7207 0 0
2
5.90125e-315 5.36716e-315
0
7 74LS251
144 1027 492 0 14 29
0 129 130 131 132 133 92 134 85 105
106 107 104 135 99
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4459 0 0
2
5.90125e-315 5.37752e-315
0
7 74LS251
144 1028 389 0 14 29
0 136 137 138 139 140 93 141 87 105
106 107 104 142 100
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3760 0 0
2
5.90125e-315 5.38788e-315
0
7 74LS251
144 1034 287 0 14 29
0 143 144 145 146 147 94 148 88 105
106 107 104 149 101
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
754 0 0
2
5.90125e-315 5.39306e-315
0
7 74LS251
144 1033 187 0 14 29
0 150 151 152 153 154 95 155 89 105
106 107 104 156 102
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9767 0 0
2
5.90125e-315 5.39824e-315
0
8 Hex Key~
166 1115 33 0 11 12
0 107 106 105 157 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
7978 0 0
2
5.90125e-315 5.40342e-315
0
7 74LS251
144 1033 94 0 14 29
0 158 159 160 161 162 78 163 78 105
106 107 104 164 103
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3142 0 0
2
5.90125e-315 5.4086e-315
0
12 Hex Display~
7 1859 45 0 18 19
10 96 97 98 99 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3284 0 0
2
5.90125e-315 5.41378e-315
0
8 Hex Key~
166 15 40 0 11 12
0 86 90 91 78 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
659 0 0
2
5.90125e-315 5.41896e-315
0
6 74136~
219 89 163 0 3 22
0 91 78 95
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3800 0 0
2
5.90125e-315 5.42414e-315
0
12 Hex Display~
7 1799 42 0 18 19
10 100 101 102 103 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6792 0 0
2
5.90125e-315 5.42933e-315
0
6 74136~
219 138 193 0 3 22
0 95 90 94
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3701 0 0
2
5.90125e-315 5.43192e-315
0
8 Hex Key~
166 52 42 0 11 12
0 5 6 7 12 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6316 0 0
2
5.90125e-315 5.43451e-315
0
233
4 0 0 0 0 0 0 74 0 0 106 2
556 1092
43 1092
3 0 0 0 0 0 0 74 0 0 104 2
556 1083
55 1083
2 4 0 0 0 0 0 74 7 0 0 4
556 1074
378 1074
378 1000
370 1000
4 1 0 0 0 0 0 8 74 0 0 4
369 927
548 927
548 1065
556 1065
1 0 5 0 0 4096 0 4 0 0 103 2
105 1009
61 1009
1 0 6 0 0 4096 0 5 0 0 104 2
148 1000
55 1000
1 0 7 0 0 4096 0 6 0 0 105 2
188 991
49 991
3 2 8 0 0 4224 0 7 4 0 0 2
325 1009
141 1009
2 2 9 0 0 4224 0 7 5 0 0 2
325 1000
184 1000
2 1 10 0 0 4224 0 6 7 0 0 2
224 991
325 991
0 3 5 0 0 4096 0 0 8 103 0 2
61 936
324 936
1 0 6 0 0 4096 0 3 0 0 104 2
168 927
55 927
2 2 11 0 0 4224 0 3 8 0 0 2
204 927
324 927
1 0 7 0 0 4096 0 8 0 0 105 2
324 918
49 918
5 7 13 0 0 8320 0 15 75 0 0 4
595 2173
626 2173
626 1970
812 1970
6 5 14 0 0 4224 0 75 23 0 0 4
812 1964
595 1964
595 1976
587 1976
5 5 15 0 0 8320 0 39 75 0 0 4
579 1776
644 1776
644 1958
812 1958
4 3 16 0 0 8320 0 75 56 0 0 4
812 1952
589 1952
589 1528
557 1528
3 5 17 0 0 8320 0 75 66 0 0 4
812 1946
636 1946
636 1320
556 1320
5 2 18 0 0 8320 0 72 75 0 0 4
601 1174
668 1174
668 1940
812 1940
1 9 2 0 0 8320 0 73 75 0 0 4
983 923
979 923
979 1955
890 1955
1 5 19 0 0 8320 0 75 74 0 0 4
812 1934
631 1934
631 1078
606 1078
8 1 20 0 0 8320 0 75 1 0 0 3
812 1976
791 1976
791 2334
1 0 7 0 0 4096 0 12 0 0 105 2
378 2250
49 2250
1 0 6 0 0 0 0 9 0 0 104 2
200 2268
55 2268
2 2 21 0 0 4224 0 9 12 0 0 2
236 2268
378 2268
2 0 6 0 0 0 0 13 0 0 104 2
321 2233
55 2233
1 0 7 0 0 0 0 10 0 0 105 2
191 2215
49 2215
2 1 22 0 0 4224 0 10 13 0 0 2
227 2215
321 2215
2 0 6 0 0 0 0 14 0 0 104 2
370 2190
55 2190
1 0 5 0 0 0 0 11 0 0 103 2
205 2172
61 2172
2 1 23 0 0 4224 0 11 14 0 0 2
241 2172
370 2172
4 3 24 0 0 12416 0 15 12 0 0 4
545 2187
516 2187
516 2259
423 2259
3 3 25 0 0 12416 0 15 13 0 0 4
545 2178
470 2178
470 2224
366 2224
3 2 26 0 0 12416 0 14 15 0 0 4
415 2181
451 2181
451 2169
545 2169
1 0 12 0 0 0 0 15 0 0 106 2
545 2160
43 2160
3 4 27 0 0 4224 0 20 23 0 0 4
392 2070
529 2070
529 1990
537 1990
3 3 28 0 0 12416 0 21 23 0 0 4
388 2018
421 2018
421 1981
537 1981
1 0 6 0 0 0 0 16 0 0 104 2
218 2079
55 2079
1 0 7 0 0 0 0 21 0 0 105 2
343 2009
49 2009
2 2 29 0 0 4224 0 16 20 0 0 2
254 2079
347 2079
1 0 7 0 0 0 0 20 0 0 105 2
347 2061
49 2061
1 0 5 0 0 0 0 17 0 0 103 2
218 2027
61 2027
2 2 30 0 0 4224 0 17 21 0 0 2
254 2027
343 2027
3 2 31 0 0 12416 0 22 23 0 0 4
330 1982
381 1982
381 1972
537 1972
2 2 32 0 0 4224 0 22 19 0 0 2
285 1991
165 1991
2 1 33 0 0 4224 0 18 22 0 0 2
222 1973
285 1973
1 0 5 0 0 0 0 19 0 0 103 2
129 1991
61 1991
1 0 6 0 0 0 0 18 0 0 104 2
186 1973
55 1973
1 0 12 0 0 0 0 23 0 0 106 2
537 1963
43 1963
5 2 34 0 0 8320 0 28 39 0 0 3
435 1784
435 1772
529 1772
1 0 5 0 0 0 0 26 0 0 103 2
258 1365
61 1365
1 0 6 0 0 0 0 25 0 0 104 2
227 1374
55 1374
1 0 12 0 0 0 0 24 0 0 106 2
199 1383
43 1383
3 2 35 0 0 4224 0 27 24 0 0 2
357 1383
235 1383
2 2 36 0 0 4224 0 25 27 0 0 2
263 1374
357 1374
2 1 37 0 0 4224 0 26 27 0 0 2
294 1365
357 1365
4 3 38 0 0 12416 0 27 66 0 0 4
402 1374
422 1374
422 1325
506 1325
1 0 7 0 0 4096 0 28 0 0 105 2
390 1771
49 1771
3 0 5 0 0 4096 0 28 0 0 103 2
390 1789
61 1789
4 2 39 0 0 4224 0 28 29 0 0 2
390 1798
215 1798
2 2 40 0 0 4224 0 33 28 0 0 2
194 1780
390 1780
1 0 12 0 0 0 0 29 0 0 106 2
179 1798
43 1798
0 1 5 0 0 0 0 0 32 103 0 2
61 1732
269 1732
0 1 7 0 0 0 0 0 31 105 0 2
49 1741
199 1741
1 0 12 0 0 0 0 30 0 0 106 2
115 1750
43 1750
2 1 41 0 0 4224 0 32 38 0 0 2
305 1732
417 1732
2 2 42 0 0 4224 0 38 31 0 0 2
417 1741
235 1741
2 3 43 0 0 4224 0 30 38 0 0 2
151 1750
417 1750
1 0 6 0 0 0 0 33 0 0 104 2
158 1780
55 1780
1 0 5 0 0 0 0 35 0 0 103 2
147 1892
61 1892
2 2 44 0 0 4224 0 35 36 0 0 2
183 1892
358 1892
1 0 12 0 0 0 0 36 0 0 106 2
358 1874
43 1874
2 0 6 0 0 0 0 37 0 0 104 2
401 1846
55 1846
2 1 45 0 0 4224 0 34 37 0 0 2
190 1828
401 1828
1 0 5 0 0 0 0 34 0 0 103 2
154 1828
61 1828
4 3 46 0 0 12416 0 39 36 0 0 4
529 1790
497 1790
497 1883
403 1883
3 3 47 0 0 12416 0 37 39 0 0 4
446 1837
464 1837
464 1781
529 1781
4 1 48 0 0 4224 0 38 39 0 0 4
462 1741
521 1741
521 1763
529 1763
1 0 5 0 0 0 0 40 0 0 103 2
127 1685
61 1685
2 3 49 0 0 4224 0 40 51 0 0 2
163 1685
341 1685
2 0 6 0 0 0 0 51 0 0 104 2
341 1676
55 1676
1 0 12 0 0 0 0 41 0 0 106 2
183 1667
43 1667
2 1 50 0 0 4224 0 41 51 0 0 2
219 1667
341 1667
1 0 7 0 0 0 0 42 0 0 105 2
152 1622
49 1622
2 2 51 0 0 4224 0 42 54 0 0 2
188 1622
299 1622
1 0 12 0 0 0 0 43 0 0 106 2
75 1613
43 1613
2 1 52 0 0 4224 0 43 54 0 0 2
111 1613
299 1613
3 0 6 0 0 0 0 54 0 0 104 2
299 1631
55 1631
4 2 53 0 0 4224 0 51 57 0 0 4
386 1676
412 1676
412 1655
420 1655
4 1 54 0 0 4224 0 54 57 0 0 4
344 1622
412 1622
412 1637
420 1637
4 3 55 0 0 8320 0 52 58 0 0 4
387 1568
402 1568
402 1515
410 1515
1 0 6 0 0 0 0 44 0 0 104 2
235 1577
55 1577
1 0 7 0 0 0 0 45 0 0 105 2
156 1568
49 1568
2 3 56 0 0 4224 0 44 52 0 0 2
271 1577
342 1577
2 2 57 0 0 4224 0 45 52 0 0 2
192 1568
342 1568
1 0 12 0 0 0 0 52 0 0 106 2
342 1559
43 1559
3 0 5 0 0 0 0 53 0 0 103 2
299 1543
61 1543
1 0 6 0 0 0 0 46 0 0 104 2
206 1534
55 1534
4 2 58 0 0 4224 0 53 58 0 0 4
344 1534
381 1534
381 1506
411 1506
2 2 59 0 0 4224 0 46 53 0 0 2
242 1534
299 1534
0 1 7 0 0 0 0 0 53 105 0 2
49 1525
299 1525
1 4 5 0 0 4224 0 110 47 0 0 2
61 66
61 2334
2 3 6 0 0 4224 0 110 47 0 0 2
55 66
55 2334
3 2 7 0 0 4224 0 110 47 0 0 2
49 66
49 2334
4 1 12 0 0 4224 0 110 47 0 0 2
43 66
43 2334
4 1 60 0 0 4224 0 55 58 0 0 2
384 1497
410 1497
2 3 61 0 0 4224 0 48 55 0 0 2
203 1506
339 1506
2 2 62 0 0 4224 0 55 49 0 0 2
339 1497
252 1497
2 1 63 0 0 4224 0 50 55 0 0 2
299 1488
339 1488
1 1 5 0 0 128 0 110 48 0 0 3
61 66
61 1506
167 1506
2 1 6 0 0 128 0 110 49 0 0 3
55 66
55 1497
216 1497
3 1 7 0 0 128 0 110 50 0 0 3
49 66
49 1488
263 1488
2 3 64 0 0 8320 0 56 57 0 0 4
511 1537
490 1537
490 1646
466 1646
4 1 65 0 0 4224 0 58 56 0 0 4
456 1506
489 1506
489 1519
511 1519
3 4 66 0 0 8320 0 59 66 0 0 4
356 1418
439 1418
439 1334
506 1334
2 2 67 0 0 4224 0 59 62 0 0 2
311 1427
186 1427
2 1 68 0 0 4224 0 63 59 0 0 2
113 1409
311 1409
2 1 6 0 0 128 0 110 62 0 0 3
55 66
55 1427
150 1427
3 1 7 0 0 128 0 110 63 0 0 3
49 66
49 1409
77 1409
4 2 69 0 0 12416 0 60 66 0 0 4
357 1342
406 1342
406 1316
506 1316
2 3 70 0 0 4224 0 64 60 0 0 2
166 1351
312 1351
1 2 6 0 0 0 0 60 110 0 0 3
312 1333
55 1333
55 66
3 2 7 0 0 0 0 110 60 0 0 3
49 66
49 1342
312 1342
4 1 12 0 0 128 0 110 64 0 0 3
43 66
43 1351
130 1351
4 1 71 0 0 4224 0 61 66 0 0 2
403 1307
506 1307
2 1 72 0 0 4224 0 65 61 0 0 2
189 1298
358 1298
4 1 12 0 0 0 0 110 65 0 0 3
43 66
43 1298
153 1298
1 2 5 0 0 0 0 110 61 0 0 3
61 66
61 1307
358 1307
2 3 6 0 0 0 0 110 61 0 0 3
55 66
55 1316
358 1316
3 4 73 0 0 12416 0 69 72 0 0 4
405 1220
471 1220
471 1188
551 1188
2 2 74 0 0 4224 0 69 67 0 0 2
360 1229
219 1229
2 1 75 0 0 4224 0 68 69 0 0 2
181 1211
360 1211
2 1 6 0 0 128 0 110 67 0 0 3
55 66
55 1229
183 1229
1 1 5 0 0 128 0 110 68 0 0 3
61 66
61 1211
145 1211
3 3 76 0 0 12416 0 70 72 0 0 4
332 1194
368 1194
368 1179
551 1179
1 2 5 0 0 0 0 110 70 0 0 3
61 66
61 1203
287 1203
2 1 6 0 0 0 0 110 70 0 0 3
55 66
55 1185
287 1185
2 2 77 0 0 4224 0 71 72 0 0 2
118 1170
551 1170
3 1 7 0 0 128 0 110 71 0 0 3
49 66
49 1170
82 1170
4 1 12 0 0 128 0 110 72 0 0 3
43 66
43 1161
551 1161
4 1 78 0 0 4096 0 106 82 0 0 3
6 64
6 439
184 439
3 8 79 0 0 4224 0 76 96 0 0 4
160 769
603 769
603 837
991 837
3 8 80 0 0 16512 0 77 97 0 0 5
162 719
162 724
577 724
577 735
995 735
3 8 81 0 0 12416 0 78 98 0 0 4
160 667
566 667
566 635
995 635
3 6 82 0 0 8320 0 91 96 0 0 4
418 355
528 355
528 819
991 819
3 6 83 0 0 12416 0 92 97 0 0 4
368 331
537 331
537 717
995 717
3 6 84 0 0 12416 0 93 98 0 0 4
317 295
550 295
550 617
995 617
1 2 5 0 0 0 0 110 76 0 0 3
61 66
61 778
111 778
2 1 6 0 0 0 0 110 76 0 0 3
55 66
55 760
111 760
2 2 6 0 0 0 0 77 110 0 0 3
113 728
55 728
55 66
3 1 7 0 0 0 0 110 77 0 0 3
49 66
49 710
113 710
3 2 7 0 0 0 0 110 78 0 0 3
49 66
49 676
111 676
4 1 12 0 0 0 0 110 78 0 0 3
43 66
43 658
111 658
3 8 85 0 0 4224 0 79 99 0 0 4
159 612
605 612
605 528
995 528
4 2 12 0 0 0 0 110 79 0 0 3
43 66
43 621
110 621
1 1 86 0 0 4224 0 106 79 0 0 3
24 64
24 603
110 603
3 8 87 0 0 4224 0 80 100 0 0 4
166 564
599 564
599 425
996 425
3 8 88 0 0 4224 0 81 101 0 0 4
159 513
592 513
592 323
1002 323
3 8 89 0 0 12416 0 82 102 0 0 4
233 448
583 448
583 223
1001 223
2 1 86 0 0 0 0 80 106 0 0 3
117 573
24 573
24 64
2 1 90 0 0 4224 0 106 80 0 0 3
18 64
18 555
117 555
2 2 90 0 0 0 0 81 106 0 0 3
110 522
18 522
18 64
3 1 91 0 0 4224 0 106 81 0 0 3
12 64
12 504
110 504
2 3 91 0 0 0 0 82 106 0 0 3
184 457
12 457
12 64
3 6 92 0 0 12416 0 94 99 0 0 4
270 266
518 266
518 510
995 510
3 6 93 0 0 12416 0 95 100 0 0 4
219 225
501 225
501 407
996 407
3 6 94 0 0 12416 0 109 101 0 0 4
171 193
511 193
511 305
1002 305
3 6 95 0 0 12416 0 107 102 0 0 4
122 163
516 163
516 205
1001 205
4 8 78 0 0 8320 0 106 104 0 0 3
6 64
6 130
1001 130
4 6 78 0 0 0 0 106 104 0 0 3
6 64
6 112
1001 112
14 1 96 0 0 8192 0 96 83 0 0 3
1055 837
1417 837
1417 52
14 1 97 0 0 8192 0 97 84 0 0 3
1059 735
1382 735
1382 42
14 1 98 0 0 8192 0 98 85 0 0 3
1059 635
1354 635
1354 41
14 1 99 0 0 8192 0 99 86 0 0 3
1059 528
1332 528
1332 41
14 1 100 0 0 8192 0 100 87 0 0 3
1060 425
1298 425
1298 45
14 1 101 0 0 8192 0 101 88 0 0 3
1066 323
1273 323
1273 49
14 1 102 0 0 4096 0 102 89 0 0 3
1065 223
1250 223
1250 51
14 1 103 0 0 4096 0 104 90 0 0 3
1065 130
1215 130
1215 52
14 1 96 0 0 4224 0 96 105 0 0 3
1055 837
1868 837
1868 69
14 2 97 0 0 4224 0 97 105 0 0 3
1059 735
1862 735
1862 69
14 3 98 0 0 4224 0 98 105 0 0 3
1059 635
1856 635
1856 69
14 4 99 0 0 4224 0 99 105 0 0 3
1059 528
1850 528
1850 69
2 1 5 0 0 0 0 91 110 0 0 3
369 364
61 364
61 66
3 1 83 0 0 0 0 92 91 0 0 4
368 331
366 331
366 346
369 346
2 2 6 0 0 0 0 92 110 0 0 3
319 340
55 340
55 66
3 1 84 0 0 0 0 93 92 0 0 3
317 295
317 322
319 322
2 3 7 0 0 0 0 93 110 0 0 3
268 304
49 304
49 66
3 1 92 0 0 0 0 94 93 0 0 3
270 266
268 266
268 286
4 2 12 0 0 0 0 110 94 0 0 3
43 66
43 275
221 275
3 1 93 0 0 0 0 95 94 0 0 4
219 225
220 225
220 257
221 257
1 2 86 0 0 0 0 106 95 0 0 3
24 64
24 234
170 234
3 1 94 0 0 0 0 109 95 0 0 4
171 193
169 193
169 216
170 216
2 2 90 0 0 0 0 106 109 0 0 3
18 64
18 202
122 202
12 1 104 0 0 8320 0 96 2 0 0 3
1061 801
1160 801
1160 34
12 1 104 0 0 0 0 97 2 0 0 3
1065 699
1160 699
1160 34
12 1 104 0 0 0 0 98 2 0 0 3
1065 599
1160 599
1160 34
12 1 104 0 0 0 0 99 2 0 0 3
1065 492
1160 492
1160 34
12 1 104 0 0 0 0 100 2 0 0 3
1066 389
1160 389
1160 34
12 1 104 0 0 0 0 101 2 0 0 3
1072 287
1160 287
1160 34
12 1 104 0 0 0 0 102 2 0 0 3
1071 187
1160 187
1160 34
1 12 104 0 0 0 0 2 104 0 0 3
1160 34
1160 94
1071 94
14 1 100 0 0 4224 0 100 108 0 0 3
1060 425
1808 425
1808 66
14 2 101 0 0 4224 0 101 108 0 0 3
1066 323
1802 323
1802 66
14 3 102 0 0 4224 0 102 108 0 0 3
1065 223
1796 223
1796 66
14 4 103 0 0 4224 0 104 108 0 0 3
1065 130
1790 130
1790 66
9 3 105 0 0 8192 0 98 103 0 0 3
1059 572
1112 572
1112 57
9 3 105 0 0 8192 0 97 103 0 0 3
1059 672
1112 672
1112 57
3 9 105 0 0 4224 0 103 96 0 0 3
1112 57
1112 774
1055 774
10 2 106 0 0 8320 0 96 103 0 0 3
1055 783
1118 783
1118 57
10 2 106 0 0 0 0 97 103 0 0 3
1059 681
1118 681
1118 57
2 10 106 0 0 0 0 103 98 0 0 3
1118 57
1118 581
1059 581
11 1 107 0 0 8320 0 96 103 0 0 3
1055 792
1124 792
1124 57
11 1 107 0 0 0 0 97 103 0 0 3
1059 690
1124 690
1124 57
11 1 107 0 0 0 0 98 103 0 0 3
1059 590
1124 590
1124 57
9 3 105 0 0 0 0 99 103 0 0 3
1059 465
1112 465
1112 57
9 3 105 0 0 0 0 100 103 0 0 3
1060 362
1112 362
1112 57
2 10 106 0 0 0 0 103 99 0 0 3
1118 57
1118 474
1059 474
2 10 106 0 0 0 0 103 100 0 0 3
1118 57
1118 371
1060 371
11 1 107 0 0 0 0 99 103 0 0 3
1059 483
1124 483
1124 57
1 11 107 0 0 0 0 103 100 0 0 3
1124 57
1124 380
1060 380
1 11 107 0 0 0 0 103 101 0 0 3
1124 57
1124 278
1066 278
10 2 106 0 0 0 0 101 103 0 0 3
1066 269
1118 269
1118 57
3 9 105 0 0 0 0 103 101 0 0 3
1112 57
1112 260
1066 260
11 1 107 0 0 0 0 102 103 0 0 3
1065 178
1124 178
1124 57
2 10 106 0 0 0 0 103 102 0 0 3
1118 57
1118 169
1065 169
9 3 105 0 0 0 0 102 103 0 0 3
1065 160
1112 160
1112 57
3 9 105 0 0 0 0 103 104 0 0 3
1112 57
1112 67
1065 67
2 10 106 0 0 0 0 103 104 0 0 3
1118 57
1118 76
1065 76
1 11 107 0 0 0 0 103 104 0 0 3
1124 57
1124 85
1065 85
3 1 91 0 0 0 0 106 107 0 0 3
12 64
12 154
73 154
4 2 78 0 0 0 0 106 107 0 0 3
6 64
6 172
73 172
3 1 95 0 0 0 0 107 109 0 0 2
122 163
122 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
