CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
176 80 1364 707
42991634 0
0
6 Title:
5 Name:
0
0
0
37
9 2-In NOR~
219 224 572 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
5130 0 0
2
45426.5 0
0
9 2-In AND~
219 394 580 0 3 22
0 6 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
391 0 0
2
45426.5 0
0
9 2-In AND~
219 238 634 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3124 0 0
2
45426.5 0
0
9 2-In AND~
219 400 410 0 3 22
0 4 10 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3421 0 0
2
45426.5 0
0
9 3-In NOR~
219 192 419 0 4 22
0 8 5 7 10
0
0 0 624 0
6 74LS27
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 6 0
1 U
8157 0 0
2
45426.5 0
0
9 2-In AND~
219 398 236 0 3 22
0 5 12 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5572 0 0
2
45426.5 0
0
9 4-In NOR~
219 264 245 0 5 22
0 8 4 7 25 12
0
0 0 624 0
4 4002
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 512 2 2 5 0
1 U
8901 0 0
2
45426.5 0
0
9 4-In NOR~
219 381 106 0 5 22
0 8 5 4 7 13
0
0 0 624 0
4 4002
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 5 0
1 U
7361 0 0
2
45426.5 0
0
9 2-In AND~
219 397 165 0 3 22
0 8 15 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4747 0 0
2
45426.5 0
0
9 3-In NOR~
219 225 174 0 4 22
0 5 4 7 15
0
0 0 624 0
6 74LS27
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
972 0 0
2
45426.5 0
0
14 Logic Display~
6 1522 55 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3472 0 0
2
45426.5 0
0
14 Logic Display~
6 1454 58 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
9998 0 0
2
45426.5 0
0
14 Logic Display~
6 1388 62 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3536 0 0
2
45426.5 0
0
14 Logic Display~
6 1331 67 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
4597 0 0
2
45426.5 0
0
14 Logic Display~
6 1261 68 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3835 0 0
2
45426.5 0
0
14 Logic Display~
6 1192 64 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3670 0 0
2
45426.5 0
0
14 Logic Display~
6 919 58 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
5616 0 0
2
45426.5 0
0
14 Logic Display~
6 841 47 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
9323 0 0
2
45426.5 0
0
14 Logic Display~
6 654 46 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
45426.5 0
0
14 Logic Display~
6 586 40 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45426.5 0
0
14 Logic Display~
6 521 44 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
45426.5 0
0
14 Logic Display~
6 486 47 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45426.5 0
0
14 Logic Display~
6 447 47 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
45426.5 0
0
9 2-In AND~
219 439 829 0 3 22
0 17 18 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6369 0 0
2
45426.5 0
0
9 2-In NOR~
219 199 893 0 3 22
0 5 4 18
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9172 0 0
2
45426.5 0
0
9 2-In AND~
219 393 486 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7100 0 0
2
45426.5 0
0
9 2-In NOR~
219 184 522 0 3 22
0 5 7 20
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3820 0 0
2
45426.5 0
0
9 2-In NOR~
219 198 290 0 3 22
0 4 7 22
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7678 0 0
2
45426.5 0
0
9 2-In AND~
219 401 299 0 3 22
0 22 24 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
961 0 0
2
45426.5 0
0
9 2-In AND~
219 212 821 0 3 22
0 8 7 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3178 0 0
2
45426.5 0
0
9 2-In AND~
219 217 477 0 3 22
0 8 4 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3409 0 0
2
45426.5 0
0
9 2-In AND~
219 204 349 0 3 22
0 8 5 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
45426.5 0
0
14 Logic Display~
6 1018 62 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
45426.5 0
0
14 Logic Display~
6 620 39 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
45426.5 0
0
12 Hex Display~
7 50 256 0 16 19
10 34 35 36 37 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
9265 0 0
2
45426.5 0
0
14 Logic Display~
6 551 39 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
45426.5 0
0
8 Hex Key~
166 110 60 0 11 12
0 8 5 4 7 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9424 0 0
2
45426.5 0
0
51
3 1 2 0 0 8320 0 2 19 0 0 3
415 580
654 580
654 64
3 2 3 0 0 12432 0 3 2 0 0 4
259 634
262 634
262 589
370 589
2 3 4 0 0 8192 0 3 37 0 0 3
214 643
107 643
107 84
2 1 5 0 0 4096 0 37 3 0 0 3
113 84
113 625
214 625
3 1 6 0 0 8320 0 1 2 0 0 3
263 572
263 571
370 571
2 4 7 0 0 8192 0 1 37 0 0 3
211 581
101 581
101 84
1 1 8 0 0 4096 0 37 1 0 0 3
119 84
119 563
211 563
3 1 9 0 0 8320 0 4 20 0 0 3
421 410
586 410
586 58
3 4 7 0 0 0 0 5 37 0 0 3
179 428
101 428
101 84
2 2 5 0 0 0 0 37 5 0 0 3
113 84
113 419
180 419
1 1 8 0 0 0 0 5 37 0 0 3
179 410
119 410
119 84
2 4 10 0 0 4224 0 4 5 0 0 2
376 419
231 419
3 1 4 0 0 0 0 37 4 0 0 3
107 84
107 401
376 401
3 1 11 0 0 8320 0 6 21 0 0 3
419 236
521 236
521 62
2 5 12 0 0 4224 0 6 7 0 0 2
374 245
303 245
2 1 5 0 0 0 0 37 6 0 0 3
113 84
113 227
374 227
3 4 7 0 0 0 0 7 37 0 0 3
247 250
101 250
101 84
3 2 4 0 0 0 0 37 7 0 0 3
107 84
107 241
247 241
1 1 8 0 0 0 0 37 7 0 0 3
119 84
119 232
247 232
5 1 13 0 0 8320 0 8 23 0 0 3
420 106
447 106
447 65
4 4 7 0 0 0 0 8 37 0 0 3
364 120
101 120
101 84
3 3 4 0 0 0 0 8 37 0 0 3
364 111
107 111
107 84
2 2 5 0 0 0 0 8 37 0 0 3
364 102
113 102
113 84
1 1 8 0 0 0 0 37 8 0 0 3
119 84
119 93
364 93
3 1 14 0 0 8320 0 9 22 0 0 3
418 165
486 165
486 65
2 4 15 0 0 4224 0 9 10 0 0 2
373 174
264 174
1 1 8 0 0 0 0 37 9 0 0 3
119 84
119 156
373 156
3 4 7 0 0 0 0 10 37 0 0 3
212 183
101 183
101 84
2 3 4 0 0 0 0 10 37 0 0 3
213 174
107 174
107 84
2 1 5 0 0 0 0 37 10 0 0 3
113 84
113 165
212 165
3 1 16 0 0 8320 0 24 33 0 0 3
460 829
1018 829
1018 80
3 1 17 0 0 4224 0 30 24 0 0 4
233 821
361 821
361 820
415 820
3 2 18 0 0 4224 0 25 24 0 0 3
238 893
415 893
415 838
3 2 4 0 0 4224 0 37 25 0 0 3
107 84
107 902
186 902
2 1 5 0 0 4224 0 37 25 0 0 3
113 84
113 884
186 884
3 1 19 0 0 8320 0 26 34 0 0 3
414 486
620 486
620 57
3 2 20 0 0 12416 0 27 26 0 0 4
223 522
254 522
254 495
369 495
3 1 21 0 0 4224 0 31 26 0 0 2
238 477
369 477
4 2 7 0 0 0 0 37 27 0 0 3
101 84
101 531
171 531
2 1 5 0 0 128 0 37 27 0 0 3
113 84
113 513
171 513
3 1 22 0 0 4224 0 28 29 0 0 2
237 290
377 290
4 2 7 0 0 0 0 37 28 0 0 3
101 84
101 299
185 299
3 1 4 0 0 0 0 37 28 0 0 3
107 84
107 281
185 281
3 1 23 0 0 8320 0 29 36 0 0 3
422 299
551 299
551 57
3 2 24 0 0 4224 0 32 29 0 0 4
225 349
311 349
311 308
377 308
4 2 7 0 0 4224 0 37 30 0 0 3
101 84
101 830
188 830
1 1 8 0 0 4224 0 37 30 0 0 3
119 84
119 812
188 812
3 2 4 0 0 128 0 37 31 0 0 3
107 84
107 486
193 486
1 1 8 0 0 0 0 37 31 0 0 3
119 84
119 468
193 468
2 2 5 0 0 128 0 37 32 0 0 3
113 84
113 358
180 358
1 1 8 0 0 0 0 37 32 0 0 3
119 84
119 340
180 340
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
