CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
470 0 1 90 10
1712 80 2814 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
2263 80 2814 659
9437202 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 1084 83 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
951 0 0
2
45075.8 0
0
13 Logic Switch~
5 257 977 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-31 -1 -17 7
2 V2
-30 -12 -16 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9536 0 0
2
45075.8 0
0
13 Logic Switch~
5 226 708 0 1 11
0 2
0
0 0 21360 0
2 0V
-30 3 -16 11
2 V1
-29 -7 -15 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5495 0 0
2
45075.8 0
0
7 74LS251
144 898 172 0 14 29
0 2 4 2 5 6 7 8 9 19
20 21 3 48 18
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8152 0 0
2
45075.9 0
0
7 74LS251
144 894 299 0 14 29
0 2 10 11 12 13 14 15 16 19
20 21 3 49 17
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U7
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
6223 0 0
2
45075.9 0
0
12 Hex Display~
7 1155 76 0 16 19
10 39 40 41 42 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5441 0 0
2
45075.8 1
0
12 Hex Display~
7 1214 75 0 18 19
10 18 17 37 38 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3189 0 0
2
45075.8 0
0
8 Hex Key~
166 1022 73 0 11 12
0 21 20 19 50 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
8460 0 0
2
45075.8 0
0
7 74LS251
144 897 1056 0 14 29
0 2 2 35 2 2 2 2 2 19
20 21 3 51 42
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U14
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
5179 0 0
2
45075.8 0
0
7 74LS251
144 896 924 0 14 29
0 2 36 33 2 2 2 2 2 19
20 21 3 52 41
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U13
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3593 0 0
2
45075.8 0
0
7 74LS251
144 894 799 0 14 29
0 2 35 28 2 2 2 2 2 19
20 21 3 53 40
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3928 0 0
2
45075.8 0
0
7 74LS251
144 895 675 0 14 29
0 2 33 22 2 2 34 2 2 19
20 21 3 54 39
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
363 0 0
2
45075.8 0
0
7 74LS251
144 894 554 0 14 29
0 2 28 10 2 29 30 31 32 19
20 21 3 55 38
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8132 0 0
2
45075.8 0
0
7 74LS251
144 895 415 0 14 29
0 2 22 4 23 24 25 26 27 19
20 21 3 56 37
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
65 0 0
2
45075.8 0
0
6 74LS85
106 319 1101 0 14 29
0 36 35 33 28 22 10 4 11 57
58 59 23 12 5
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
6609 0 0
2
45075.8 0
0
9 Inverter~
13 251 834 0 2 22
0 22 44
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
8995 0 0
2
45075.8 3
0
9 Inverter~
13 251 871 0 2 22
0 10 45
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3918 0 0
2
45075.8 2
0
9 Inverter~
13 251 942 0 2 22
0 11 47
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
7519 0 0
2
45075.8 1
0
9 Inverter~
13 251 906 0 2 22
0 4 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
377 0 0
2
45075.8 0
0
4 4008
219 389 891 0 14 29
0 36 35 33 28 44 45 46 47 43
6 13 24 29 60
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
8816 0 0
2
45075.8 0
0
4 4008
219 417 661 0 14 29
0 36 35 33 28 22 10 4 11 2
7 14 25 30 34
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 0 0 0 0
1 U
3877 0 0
2
45075.8 0
0
9 2-In AND~
219 257 531 0 3 22
0 22 36 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
926 0 0
2
45075.8 0
0
9 2-In AND~
219 258 482 0 3 22
0 10 35 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7262 0 0
2
45075.8 0
0
9 2-In AND~
219 258 429 0 3 22
0 4 33 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5267 0 0
2
45075.8 0
0
9 2-In AND~
219 259 376 0 3 22
0 11 28 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8838 0 0
2
45075.8 0
0
8 2-In OR~
219 251 320 0 3 22
0 22 36 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7159 0 0
2
45075.8 0
0
8 2-In OR~
219 253 268 0 3 22
0 10 35 27
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5812 0 0
2
45075.8 0
0
8 2-In OR~
219 254 213 0 3 22
0 4 33 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
331 0 0
2
45075.8 0
0
8 2-In OR~
219 254 157 0 3 22
0 11 28 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9604 0 0
2
45075.8 0
0
8 Hex Key~
166 108 57 0 11 12
0 28 33 35 36 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7518 0 0
2
45075.8 0
0
8 Hex Key~
166 163 58 0 11 12
0 11 4 10 22 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4832 0 0
2
45075.8 0
0
150
1 8 2 0 0 8336 0 3 12 0 0 5
238 708
238 729
756 729
756 711
863 711
1 1 2 0 0 0 0 4 5 0 0 4
866 145
830 145
830 272
862 272
1 12 3 0 0 8192 0 1 4 0 0 3
1084 95
1084 172
936 172
1 4 2 0 0 0 0 13 13 0 0 4
862 527
854 527
854 554
862 554
2 2 4 0 0 4096 0 4 31 0 0 5
866 154
364 154
364 122
166 122
166 82
1 3 2 0 0 0 0 4 4 0 0 4
866 145
804 145
804 163
866 163
4 14 5 0 0 8320 0 4 15 0 0 4
866 172
685 172
685 1137
351 1137
5 10 6 0 0 8320 0 4 20 0 0 4
866 181
655 181
655 900
421 900
6 10 7 0 0 8320 0 4 21 0 0 4
866 190
591 190
591 670
449 670
3 7 8 0 0 4224 0 25 4 0 0 4
280 376
780 376
780 199
866 199
3 8 9 0 0 12416 0 29 4 0 0 4
287 157
312 157
312 208
866 208
2 3 10 0 0 4096 0 5 31 0 0 5
862 281
451 281
451 109
160 109
160 82
3 1 11 0 0 12288 0 5 31 0 0 4
862 290
560 290
560 82
172 82
4 13 12 0 0 8320 0 5 15 0 0 4
862 299
629 299
629 1128
351 1128
11 5 13 0 0 8320 0 20 5 0 0 4
421 891
616 891
616 308
862 308
6 11 14 0 0 4224 0 5 21 0 0 4
862 317
469 317
469 661
449 661
3 7 15 0 0 12416 0 24 5 0 0 4
279 429
433 429
433 326
862 326
8 3 16 0 0 4224 0 5 28 0 0 6
862 335
498 335
498 252
295 252
295 213
287 213
12 1 3 0 0 8192 0 5 1 0 0 3
932 299
1084 299
1084 95
14 2 17 0 0 4224 0 5 7 0 0 3
926 335
1217 335
1217 99
14 1 18 0 0 4224 0 4 7 0 0 3
930 208
1223 208
1223 99
3 9 19 0 0 4096 0 8 5 0 0 3
1019 97
1019 272
926 272
2 10 20 0 0 4096 0 8 5 0 0 3
1025 97
1025 281
926 281
1 11 21 0 0 4096 0 8 5 0 0 3
1031 97
1031 290
926 290
3 9 19 0 0 0 0 8 4 0 0 3
1019 97
1019 145
930 145
2 10 20 0 0 0 0 8 4 0 0 3
1025 97
1025 154
930 154
1 11 21 0 0 0 0 8 4 0 0 3
1031 97
1031 163
930 163
1 1 2 0 0 0 0 5 14 0 0 4
862 272
791 272
791 388
863 388
2 4 22 0 0 4096 0 14 31 0 0 3
863 397
154 397
154 82
3 2 4 0 0 0 0 14 31 0 0 5
863 406
406 406
406 93
166 93
166 82
4 12 23 0 0 8320 0 14 15 0 0 4
863 415
563 415
563 1119
351 1119
5 12 24 0 0 8320 0 14 20 0 0 4
863 424
545 424
545 882
421 882
6 12 25 0 0 4224 0 14 21 0 0 4
863 433
482 433
482 652
449 652
3 7 26 0 0 12416 0 23 14 0 0 4
279 482
322 482
322 442
863 442
3 8 27 0 0 12416 0 27 14 0 0 4
286 268
343 268
343 451
863 451
2 4 28 0 0 4096 0 13 21 0 0 4
862 536
327 536
327 652
385 652
3 3 10 0 0 16384 0 13 31 0 0 5
862 545
386 545
386 581
160 581
160 82
13 5 29 0 0 12416 0 20 13 0 0 4
421 873
521 873
521 563
862 563
13 6 30 0 0 12416 0 21 13 0 0 4
449 643
642 643
642 572
862 572
3 7 31 0 0 20608 0 22 13 0 0 6
278 531
299 531
299 518
504 518
504 581
862 581
3 8 32 0 0 20608 0 26 13 0 0 6
284 320
312 320
312 293
456 293
456 590
862 590
1 1 2 0 0 0 0 14 13 0 0 4
863 388
729 388
729 527
862 527
1 1 2 0 0 128 0 13 12 0 0 4
862 527
700 527
700 648
863 648
2 3 33 0 0 4096 0 12 21 0 0 6
863 657
576 657
576 721
375 721
375 643
385 643
1 4 2 0 0 0 0 12 12 0 0 4
863 648
804 648
804 675
863 675
4 5 2 0 0 0 0 12 12 0 0 2
863 675
863 684
3 4 22 0 0 0 0 12 31 0 0 5
863 666
603 666
603 734
154 734
154 82
14 6 34 0 0 4224 0 21 12 0 0 5
449 625
673 625
673 692
863 692
863 693
7 5 2 0 0 0 0 12 12 0 0 4
863 702
804 702
804 684
863 684
7 8 2 0 0 0 0 12 12 0 0 2
863 702
863 711
8 8 2 0 0 0 0 12 11 0 0 4
863 711
803 711
803 835
862 835
2 2 35 0 0 12288 0 21 11 0 0 4
385 634
351 634
351 781
862 781
4 3 28 0 0 0 0 15 11 0 0 6
287 1101
250 1101
250 1162
641 1162
641 790
862 790
7 8 2 0 0 0 0 11 11 0 0 2
862 826
862 835
6 7 2 0 0 0 0 11 11 0 0 2
862 817
862 826
5 6 2 0 0 0 0 11 11 0 0 2
862 808
862 817
4 5 2 0 0 0 0 11 11 0 0 2
862 799
862 808
1 4 2 0 0 0 0 11 11 0 0 4
862 772
765 772
765 799
862 799
1 2 36 0 0 12288 0 21 10 0 0 6
385 625
299 625
299 755
669 755
669 906
864 906
3 3 33 0 0 12288 0 15 10 0 0 6
287 1092
234 1092
234 1174
669 1174
669 915
864 915
8 8 2 0 0 0 0 10 11 0 0 4
864 960
764 960
764 835
862 835
7 8 2 0 0 0 0 10 10 0 0 2
864 951
864 960
6 7 2 0 0 0 0 10 10 0 0 2
864 942
864 951
5 6 2 0 0 0 0 10 10 0 0 2
864 933
864 942
4 5 2 0 0 0 0 10 10 0 0 2
864 924
864 933
1 4 2 0 0 0 0 10 10 0 0 4
864 897
811 897
811 924
864 924
1 4 2 0 0 0 0 9 9 0 0 4
865 1029
832 1029
832 1056
865 1056
8 8 2 0 0 0 0 9 10 0 0 4
865 1092
730 1092
730 960
864 960
7 8 2 0 0 0 0 9 9 0 0 2
865 1083
865 1092
6 7 2 0 0 0 0 9 9 0 0 2
865 1074
865 1083
5 6 2 0 0 0 0 9 9 0 0 2
865 1065
865 1074
4 5 2 0 0 0 0 9 9 0 0 2
865 1056
865 1065
1 2 2 0 0 0 0 9 9 0 0 2
865 1029
865 1038
2 3 35 0 0 0 0 15 9 0 0 6
287 1083
222 1083
222 1188
692 1188
692 1047
865 1047
3 14 37 0 0 4224 0 7 14 0 0 3
1211 99
1211 451
927 451
4 14 38 0 0 4224 0 7 13 0 0 3
1205 99
1205 590
926 590
1 14 39 0 0 4224 0 6 12 0 0 3
1164 100
1164 711
927 711
2 14 40 0 0 4224 0 6 11 0 0 3
1158 100
1158 835
926 835
3 14 41 0 0 4224 0 6 10 0 0 3
1152 100
1152 960
928 960
4 14 42 0 0 4224 0 6 9 0 0 3
1146 100
1146 1092
929 1092
1 12 3 0 0 4224 0 1 9 0 0 3
1084 95
1084 1056
935 1056
1 12 3 0 0 0 0 1 10 0 0 3
1084 95
1084 924
934 924
1 12 3 0 0 0 0 1 11 0 0 3
1084 95
1084 799
932 799
1 12 3 0 0 0 0 1 12 0 0 3
1084 95
1084 675
933 675
1 12 3 0 0 0 0 1 13 0 0 3
1084 95
1084 554
932 554
1 12 3 0 0 0 0 1 14 0 0 3
1084 95
1084 415
933 415
3 9 19 0 0 4224 0 8 9 0 0 3
1019 97
1019 1029
929 1029
2 10 20 0 0 4224 0 8 9 0 0 3
1025 97
1025 1038
929 1038
1 11 21 0 0 4224 0 8 9 0 0 3
1031 97
1031 1047
929 1047
3 9 19 0 0 0 0 8 10 0 0 3
1019 97
1019 897
928 897
2 10 20 0 0 0 0 8 10 0 0 3
1025 97
1025 906
928 906
1 11 21 0 0 0 0 8 10 0 0 3
1031 97
1031 915
928 915
3 9 19 0 0 0 0 8 11 0 0 3
1019 97
1019 772
926 772
2 10 20 0 0 0 0 8 11 0 0 3
1025 97
1025 781
926 781
1 11 21 0 0 0 0 8 11 0 0 3
1031 97
1031 790
926 790
3 9 19 0 0 0 0 8 12 0 0 3
1019 97
1019 648
927 648
2 10 20 0 0 0 0 8 12 0 0 3
1025 97
1025 657
927 657
1 11 21 0 0 0 0 8 12 0 0 3
1031 97
1031 666
927 666
3 9 19 0 0 0 0 8 13 0 0 3
1019 97
1019 527
926 527
2 10 20 0 0 0 0 8 13 0 0 3
1025 97
1025 536
926 536
1 11 21 0 0 0 0 8 13 0 0 3
1031 97
1031 545
926 545
3 9 19 0 0 0 0 8 14 0 0 3
1019 97
1019 388
927 388
2 10 20 0 0 0 0 8 14 0 0 3
1025 97
1025 397
927 397
1 11 21 0 0 0 0 8 14 0 0 3
1031 97
1031 406
927 406
4 1 36 0 0 4224 0 30 15 0 0 3
99 81
99 1074
287 1074
3 2 35 0 0 4224 0 30 15 0 0 3
105 81
105 1083
287 1083
2 3 33 0 0 4224 0 30 15 0 0 3
111 81
111 1092
287 1092
1 4 28 0 0 4224 0 30 15 0 0 3
117 81
117 1101
287 1101
4 5 22 0 0 4224 0 31 15 0 0 3
154 82
154 1110
287 1110
3 6 10 0 0 4224 0 31 15 0 0 3
160 82
160 1119
287 1119
2 7 4 0 0 4224 0 31 15 0 0 3
166 82
166 1128
287 1128
1 8 11 0 0 4224 0 31 15 0 0 3
172 82
172 1137
287 1137
1 9 43 0 0 12416 0 2 20 0 0 4
269 977
289 977
289 927
357 927
4 1 36 0 0 0 0 30 20 0 0 5
99 81
99 765
337 765
337 855
357 855
3 2 35 0 0 0 0 30 20 0 0 5
105 81
105 779
325 779
325 864
357 864
2 3 33 0 0 0 0 30 20 0 0 5
111 81
111 793
315 793
315 873
357 873
1 4 28 0 0 0 0 30 20 0 0 5
117 81
117 807
301 807
301 882
357 882
4 1 22 0 0 0 0 31 16 0 0 3
154 82
154 834
236 834
3 1 10 0 0 0 0 31 17 0 0 3
160 82
160 871
236 871
2 1 4 0 0 0 0 31 19 0 0 3
166 82
166 906
236 906
1 1 11 0 0 0 0 31 18 0 0 3
172 82
172 942
236 942
2 5 44 0 0 12416 0 16 20 0 0 4
272 834
289 834
289 891
357 891
2 6 45 0 0 12416 0 17 20 0 0 4
272 871
280 871
280 900
357 900
2 7 46 0 0 8320 0 19 20 0 0 3
272 906
272 909
357 909
2 8 47 0 0 12416 0 18 20 0 0 4
272 942
280 942
280 918
357 918
4 1 36 0 0 0 0 30 21 0 0 3
99 81
99 625
385 625
3 2 35 0 0 0 0 30 21 0 0 3
105 81
105 634
385 634
2 3 33 0 0 0 0 30 21 0 0 3
111 81
111 643
385 643
1 4 28 0 0 0 0 30 21 0 0 3
117 81
117 652
385 652
4 5 22 0 0 0 0 31 21 0 0 3
154 82
154 661
385 661
3 6 10 0 0 0 0 31 21 0 0 3
160 82
160 670
385 670
2 7 4 0 0 0 0 31 21 0 0 3
166 82
166 679
385 679
1 8 11 0 0 0 0 31 21 0 0 3
172 82
172 688
385 688
1 9 2 0 0 128 0 3 21 0 0 4
238 708
264 708
264 697
385 697
4 2 36 0 0 0 0 30 22 0 0 3
99 81
99 540
233 540
3 2 35 0 0 0 0 30 23 0 0 3
105 81
105 491
234 491
2 2 33 0 0 0 0 30 24 0 0 3
111 81
111 438
234 438
1 2 28 0 0 0 0 30 25 0 0 3
117 81
117 385
235 385
4 2 36 0 0 0 0 30 26 0 0 3
99 81
99 329
238 329
3 2 35 0 0 0 0 30 27 0 0 3
105 81
105 277
240 277
2 2 33 0 0 0 0 30 28 0 0 3
111 81
111 222
241 222
1 2 28 0 0 0 0 30 29 0 0 3
117 81
117 166
241 166
4 1 22 0 0 0 0 31 22 0 0 3
154 82
154 522
233 522
3 1 10 0 0 0 0 31 23 0 0 3
160 82
160 473
234 473
2 1 4 0 0 0 0 31 24 0 0 3
166 82
166 420
234 420
1 1 11 0 0 0 0 31 25 0 0 3
172 82
172 367
235 367
4 1 22 0 0 0 0 31 26 0 0 3
154 82
154 311
238 311
3 1 10 0 0 0 0 31 27 0 0 3
160 82
160 259
240 259
2 1 4 0 0 0 0 31 28 0 0 3
166 82
166 204
241 204
1 1 11 0 0 0 0 31 29 0 0 3
172 82
172 148
241 148
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1275 75 1334 99
1286 84 1322 100
6 1= A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1274 55 1333 79
1285 64 1321 80
6 2= A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1276 37 1335 61
1287 46 1323 62
6 4= B>A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
296 1010 341 1034
306 1018 330 1034
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
366 801 411 825
376 809 400 825
3 A-B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
395 575 440 599
405 583 429 599
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
150 -3 179 21
160 5 168 21
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
95 -2 124 22
105 6 113 22
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
