CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 221 75 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
513 0 0
2
44902.5 0
0
13 Logic Switch~
5 156 274 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5737 0 0
2
44902.5 0
0
14 Logic Display~
6 356 91 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9982 0 0
2
44902.5 0
0
14 Logic Display~
6 472 170 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9576 0 0
2
44902.5 0
0
6 JK RN~
219 399 220 0 6 22
0 5 2 5 6 7 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
3507 0 0
2
44902.5 0
0
6 JK RN~
219 284 136 0 6 22
0 3 2 3 6 8 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3494 0 0
2
44902.5 0
0
9 Data Seq~
170 99 112 0 17 21
0 9 10 11 12 13 14 15 2 16
17 15 1 20 1 1 0 33
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
21 type:source { TW=100}
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
7897 0 0
2
44902.5 0
0
AAAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAAAAAAAAAAAAAAAAAAAAAAA
10
8 2 2 0 0 4096 0 7 6 0 0 4
131 148
245 148
245 128
253 128
1 3 3 0 0 4096 0 6 6 0 0 4
260 119
235 119
235 137
260 137
1 1 3 0 0 8320 0 1 6 0 0 3
221 87
221 119
260 119
6 1 4 0 0 4224 0 5 4 0 0 3
423 203
472 203
472 188
1 3 5 0 0 4096 0 5 5 0 0 4
375 203
355 203
355 221
375 221
6 1 5 0 0 8320 0 6 5 0 0 4
308 119
360 119
360 203
375 203
6 1 5 0 0 0 0 6 3 0 0 3
308 119
356 119
356 109
4 4 6 0 0 8192 0 5 6 0 0 6
399 251
399 266
283 266
283 175
284 175
284 167
4 1 6 0 0 8320 0 5 2 0 0 3
399 251
399 274
168 274
2 2 2 0 0 12432 0 6 5 0 0 4
253 128
241 128
241 212
368 212
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
4.83693e-315 0 5.23039e-315 1.58404e-314 4.83693e-315 4.83693e-315
16 0
0 0.0002 10
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
4.80864e-315 0 5.27183e-315 1.58818e-314 4.80864e-315 5.31328e-315
16 0
0 5e-06 10
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
5.7175e-315 5.26354e-315 5.31304e-315 0 5.71746e-315 5.71746e-315
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
6.08861e-315 5.26354e-315 1.38842e-314 0 6.08861e-315 6.08861e-315
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
