CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
350 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
167
13 Logic Switch~
5 1732 151 0 1 11
0 9
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90125e-315 0
0
13 Logic Switch~
5 1160 22 0 1 11
0 17
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90125e-315 5.26354e-315
0
9 CC 7-Seg~
183 1540 86 0 15 19
10 16 15 14 13 12 11 10 9 2
1 1 1 1 1 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.90125e-315 0
0
7 74LS251
144 1042 1453 0 14 29
0 166 167 168 169 170 171 18 172 6
7 8 17 173 10
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U58
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3421 0 0
2
5.90125e-315 0
0
7 74LS251
144 1039 1355 0 14 29
0 174 175 176 177 178 179 19 180 6
7 8 17 181 11
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U57
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8157 0 0
2
5.90125e-315 0
0
7 74LS251
144 1036 1250 0 14 29
0 182 183 184 185 186 187 20 188 6
7 8 17 189 12
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U56
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
5.90125e-315 0
0
7 74LS251
144 1033 1140 0 14 29
0 190 191 192 193 194 195 25 196 6
7 8 17 197 13
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U55
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8901 0 0
2
5.90125e-315 0
0
7 74LS251
144 1032 1025 0 14 29
0 198 199 200 201 202 203 26 204 6
7 8 17 205 14
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U54
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.90125e-315 0
0
7 74LS251
144 1026 921 0 14 29
0 206 207 208 209 210 211 27 212 6
7 8 17 213 15
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U53
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.90125e-315 0
0
7 Buffer~
58 950 1880 0 2 22
0 30 19
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U52B
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 47 0
1 U
972 0 0
2
5.90125e-315 0
0
7 Buffer~
58 984 1908 0 2 22
0 29 18
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U52A
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 47 0
1 U
3472 0 0
2
5.90125e-315 0
0
7 Buffer~
58 900 1349 0 2 22
0 21 25
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42F
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 37 0
1 U
9998 0 0
2
5.90125e-315 0
0
7 Buffer~
58 881 1225 0 2 22
0 22 26
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42E
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 5 37 0
1 U
3536 0 0
2
5.90125e-315 0
0
7 Buffer~
58 856 1221 0 2 22
0 23 27
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42D
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 37 0
1 U
4597 0 0
2
5.90125e-315 0
0
7 Buffer~
58 824 1223 0 2 22
0 24 28
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42C
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 37 0
1 U
3835 0 0
2
5.90125e-315 0
0
9 Inverter~
13 264 3403 0 2 22
0 4 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U49D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 44 0
1 U
3670 0 0
2
5.90125e-315 0
0
9 Inverter~
13 150 3345 0 2 22
0 3 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U49C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 44 0
1 U
5616 0 0
2
5.90125e-315 0
0
9 Inverter~
13 200 3316 0 2 22
0 36 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U49B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 44 0
1 U
9323 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 517 3394 0 3 22
0 3 34 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U51B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 46 0
1 U
317 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 418 3354 0 3 22
0 35 4 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U51A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 46 0
1 U
3108 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 345 3307 0 3 22
0 4 37 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 43 0
1 U
4299 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 785 3294 0 5 22
0 5 33 31 32 29
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U50A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 45 0
1 U
9672 0 0
2
5.90125e-315 0
0
9 Inverter~
13 184 3253 0 2 22
0 4 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U49A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 44 0
1 U
7876 0 0
2
5.90125e-315 0
0
9 Inverter~
13 232 3207 0 2 22
0 36 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 42 0
1 U
6369 0 0
2
5.90125e-315 0
0
9 Inverter~
13 235 3162 0 2 22
0 36 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 42 0
1 U
9172 0 0
2
5.90125e-315 0
0
9 Inverter~
13 197 3144 0 2 22
0 4 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 42 0
1 U
7100 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 466 3244 0 3 22
0 3 38 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 43 0
1 U
3820 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 424 3198 0 3 22
0 3 39 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 43 0
1 U
7678 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 390 3153 0 3 22
0 41 40 44
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 43 0
1 U
961 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 716 3134 0 5 22
0 5 44 43 42 30
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U40B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 35 0
1 U
3178 0 0
2
5.90125e-315 0
0
9 Inverter~
13 148 3090 0 2 22
0 36 45
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 42 0
1 U
3409 0 0
2
5.90125e-315 0
0
9 Inverter~
13 130 3040 0 2 22
0 36 46
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 42 0
1 U
3951 0 0
2
5.90125e-315 0
0
9 Inverter~
13 216 3031 0 2 22
0 4 47
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U47A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 42 0
1 U
8885 0 0
2
5.90125e-315 0
0
9 Inverter~
13 297 3022 0 2 22
0 3 48
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 40 0
1 U
3780 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 381 3081 0 3 22
0 4 45 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U37D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
9265 0 0
2
5.90125e-315 0
0
5 7415~
219 380 3031 0 4 22
0 48 47 46 50
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U46A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 41 0
1 U
9442 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 727 3053 0 3 22
0 50 49 51
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U44B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 39 0
1 U
9424 0 0
2
5.90125e-315 0
0
7 Buffer~
58 924 1848 0 2 22
0 51 20
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42B
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 37 0
1 U
9968 0 0
2
5.90125e-315 0
0
9 Inverter~
13 140 2967 0 2 22
0 36 53
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 40 0
1 U
9281 0 0
2
5.90125e-315 0
0
9 Inverter~
13 237 2949 0 2 22
0 5 52
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 40 0
1 U
8464 0 0
2
5.90125e-315 0
0
9 Inverter~
13 154 2909 0 2 22
0 3 54
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 40 0
1 U
7168 0 0
2
5.90125e-315 0
0
9 Inverter~
13 214 2900 0 2 22
0 5 55
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 40 0
1 U
3171 0 0
2
5.90125e-315 0
0
9 Inverter~
13 267 2865 0 2 22
0 4 57
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U45A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 40 0
1 U
4139 0 0
2
5.90125e-315 0
0
9 Inverter~
13 193 2856 0 2 22
0 3 56
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 36 0
1 U
6435 0 0
2
5.90125e-315 0
0
9 Inverter~
13 147 2804 0 2 22
0 4 58
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 36 0
1 U
5283 0 0
2
5.90125e-315 0
0
9 Inverter~
13 185 2762 0 2 22
0 36 66
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 36 0
1 U
6874 0 0
2
5.90125e-315 0
0
9 Inverter~
13 55 2753 0 2 22
0 4 67
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 36 0
1 U
5305 0 0
2
5.90125e-315 0
0
9 Inverter~
13 97 2744 0 2 22
0 3 68
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 36 0
1 U
34 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 729 2843 0 3 22
0 59 60 69
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U44A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 39 0
1 U
969 0 0
2
5.90125e-315 0
0
5 7415~
219 383 2958 0 4 22
0 52 4 53 61
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 38 0
1 U
8402 0 0
2
5.90125e-315 0
0
5 7415~
219 382 2909 0 4 22
0 55 54 4 62
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 38 0
1 U
3751 0 0
2
5.90125e-315 0
0
5 7415~
219 381 2856 0 4 22
0 5 56 57 63
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 38 0
1 U
4292 0 0
2
5.90125e-315 0
0
5 7415~
219 319 2804 0 4 22
0 3 58 36 64
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U38C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 33 0
1 U
6118 0 0
2
5.90125e-315 0
0
5 7415~
219 317 2753 0 4 22
0 68 67 66 65
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U38B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 33 0
1 U
34 0 0
2
5.90125e-315 0
0
8 3-In OR~
219 577 2884 0 4 22
0 63 62 61 60
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U22B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 17 0
1 U
6357 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 573 2786 0 3 22
0 65 64 59
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
319 0 0
2
5.90125e-315 0
0
7 Buffer~
58 900 1811 0 2 22
0 69 21
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U42A
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 37 0
1 U
3976 0 0
2
5.90125e-315 0
0
9 Inverter~
13 212 2689 0 2 22
0 4 71
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U41A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 36 0
1 U
7634 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 574 2684 0 5 22
0 5 3 71 36 70
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U40A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 35 0
1 U
523 0 0
2
5.90125e-315 0
0
7 Buffer~
58 881 1772 0 2 22
0 70 22
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35F
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 30 0
1 U
6748 0 0
2
5.90125e-315 0
0
9 Inverter~
13 127 2628 0 2 22
0 36 75
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 34 0
1 U
6901 0 0
2
5.90125e-315 0
0
9 Inverter~
13 175 2610 0 2 22
0 4 76
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 34 0
1 U
842 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 286 2619 0 3 22
0 76 75 73
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U37C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
3277 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 349 2573 0 3 22
0 4 36 74
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U37B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
4212 0 0
2
5.90125e-315 0
0
9 Inverter~
13 135 2550 0 2 22
0 3 77
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 34 0
1 U
4720 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 561 2554 0 5 22
0 5 77 74 73 72
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U36B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 31 0
1 U
5551 0 0
2
5.90125e-315 0
0
7 Buffer~
58 856 1759 0 2 22
0 72 23
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35E
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 5 30 0
1 U
6986 0 0
2
5.90125e-315 0
0
7 Buffer~
58 824 1765 0 2 22
0 78 24
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35D
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 30 0
1 U
8745 0 0
2
5.90125e-315 0
0
9 Inverter~
13 189 2470 0 2 22
0 36 82
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 34 0
1 U
9592 0 0
2
5.90125e-315 0
0
9 Inverter~
13 105 2461 0 2 22
0 4 81
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 34 0
1 U
8748 0 0
2
5.90125e-315 0
0
9 Inverter~
13 154 2452 0 2 22
0 3 80
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U39A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 34 0
1 U
7168 0 0
2
5.90125e-315 0
0
5 7415~
219 361 2461 0 4 22
0 80 81 82 79
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U38A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 33 0
1 U
631 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 267 2420 0 3 22
0 3 36 83
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U37A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
9466 0 0
2
5.90125e-315 0
0
8 4-In OR~
219 556 2397 0 5 22
0 5 4 83 79 78
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U36A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 31 0
1 U
3266 0 0
2
5.90125e-315 0
0
7 Buffer~
58 787 1222 0 2 22
0 87 84
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35C
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 30 0
1 U
7693 0 0
2
5.90125e-315 0
0
7 Buffer~
58 758 1220 0 2 22
0 88 85
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35B
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 30 0
1 U
3723 0 0
2
5.90125e-315 0
0
7 Buffer~
58 726 1217 0 2 22
0 89 86
0
0 0 624 90
4 4050
-14 -19 14 -11
4 U35A
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 30 0
1 U
3440 0 0
2
5.90125e-315 0
0
7 Ground~
168 1596 12 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6263 0 0
2
5.90125e-315 0
0
9 CC 7-Seg~
183 1653 91 0 15 19
10 98 97 96 95 94 93 92 9 2
1 1 1 1 1 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
4900 0 0
2
5.90125e-315 0
0
9 Inverter~
13 129 1840 0 2 22
0 101 102
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U29A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 24 0
1 U
8783 0 0
2
5.90125e-315 0
0
9 Inverter~
13 210 1741 0 2 22
0 103 105
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U27A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
3221 0 0
2
5.90125e-315 0
0
9 Inverter~
13 157 1750 0 2 22
0 104 106
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U21A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
3215 0 0
2
5.90125e-315 0
0
9 Inverter~
13 110 1759 0 2 22
0 101 107
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 29 0
1 U
7903 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 215 1831 0 3 22
0 104 102 109
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
7121 0 0
2
5.90125e-315 0
0
5 7415~
219 273 1750 0 4 22
0 105 106 107 108
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 12 0
1 U
4484 0 0
2
5.90125e-315 0
0
8 2-In OR~
219 533 1759 0 3 22
0 108 109 89
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
5996 0 0
2
5.90125e-315 0
0
9 Inverter~
13 203 1325 0 2 22
0 104 110
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 29 0
1 U
7804 0 0
2
5.90125e-315 0
0
9 2-In AND~
219 326 947 0 3 22
0 101 103 112
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
5523 0 0
2
5.90125e-315 0
0
9 Inverter~
13 120 1009 0 2 22
0 101 114
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 29 0
1 U
3330 0 0
2
45439.4 0
0
9 Inverter~
13 163 1000 0 2 22
0 104 115
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 29 0
1 U
3465 0 0
2
45439.4 1
0
9 Inverter~
13 203 991 0 2 22
0 103 116
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U34A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 29 0
1 U
8396 0 0
2
45439.4 2
0
5 7415~
219 349 1000 0 4 22
0 116 115 114 113
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 8 0
1 U
3685 0 0
2
45439.4 3
0
9 Inverter~
13 215 2268 0 2 22
0 104 117
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 27 0
1 U
7849 0 0
2
45439.4 4
0
9 Inverter~
13 206 2215 0 2 22
0 103 118
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 27 0
1 U
6343 0 0
2
45439.4 5
0
9 Inverter~
13 220 2172 0 2 22
0 101 119
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 27 0
1 U
7376 0 0
2
45439.4 6
0
9 2-In AND~
219 402 2259 0 3 22
0 103 117 120
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
9156 0 0
2
45439.4 7
0
9 2-In AND~
219 345 2224 0 3 22
0 118 104 121
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
5776 0 0
2
45439.4 8
0
9 2-In AND~
219 394 2181 0 3 22
0 119 104 122
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
7207 0 0
2
45439.4 9
0
8 4-In OR~
219 562 2173 0 5 22
0 111 122 121 120 87
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 25 0
1 U
4459 0 0
2
45439.4 10
0
9 Inverter~
13 233 2079 0 2 22
0 104 125
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 27 0
1 U
3760 0 0
2
45439.4 11
0
9 Inverter~
13 233 2027 0 2 22
0 101 126
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 27 0
1 U
754 0 0
2
45439.4 12
0
9 Inverter~
13 201 1973 0 2 22
0 104 129
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U32A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 27 0
1 U
9767 0 0
2
45439.4 13
0
9 Inverter~
13 144 1991 0 2 22
0 101 128
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U28F
-14 -18 14 -10
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 23 0
1 U
7978 0 0
2
45439.4 14
0
9 2-In AND~
219 371 2070 0 3 22
0 103 125 123
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
3142 0 0
2
45439.4 15
0
9 2-In AND~
219 367 2018 0 3 22
0 103 126 124
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
3284 0 0
2
45439.4 16
0
9 2-In AND~
219 309 1982 0 3 22
0 129 128 127
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U31A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
659 0 0
2
45439.4 17
0
8 4-In OR~
219 554 1976 0 5 22
0 111 127 124 123 88
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U30A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 25 0
1 U
3800 0 0
2
45439.4 18
0
9 Inverter~
13 142 1685 0 2 22
0 101 130
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 21 0
1 U
6792 0 0
2
45439.4 19
0
9 Inverter~
13 198 1667 0 2 22
0 111 131
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 20 0
1 U
3701 0 0
2
45439.4 20
0
9 Inverter~
13 167 1622 0 2 22
0 103 132
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 20 0
1 U
6316 0 0
2
45439.4 21
0
9 Inverter~
13 90 1613 0 2 22
0 111 133
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 20 0
1 U
8734 0 0
2
45439.4 22
0
9 Inverter~
13 250 1577 0 2 22
0 104 137
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 20 0
1 U
7988 0 0
2
45439.4 23
0
9 Inverter~
13 171 1568 0 2 22
0 103 138
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 20 0
1 U
3217 0 0
2
45439.4 24
0
9 Inverter~
13 221 1534 0 2 22
0 104 140
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U25A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 20 0
1 U
3965 0 0
2
45439.4 25
0
8 Hex Key~
166 55 2304 0 11 12
0 111 103 104 101 0 0 0 0 0
2 50
0
0 0 4656 180
0
4 KPD4
20 -2 48 6
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8239 0 0
2
45439.4 26
0
9 Inverter~
13 182 1506 0 2 22
0 101 142
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 14 0
1 U
828 0 0
2
45439.4 27
0
9 Inverter~
13 231 1497 0 2 22
0 104 143
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 14 0
1 U
6187 0 0
2
45439.4 28
0
9 Inverter~
13 278 1488 0 2 22
0 103 144
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 14 0
1 U
7107 0 0
2
45439.4 29
0
5 7415~
219 365 1676 0 4 22
0 131 104 130 134
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 19 0
1 U
6433 0 0
2
45439.4 30
0
5 7415~
219 366 1568 0 4 22
0 111 138 137 136
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 19 0
1 U
8559 0 0
2
45439.4 31
0
5 7415~
219 323 1534 0 4 22
0 103 140 101 139
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 19 0
1 U
3674 0 0
2
45439.4 32
0
5 7415~
219 323 1622 0 4 22
0 133 132 104 135
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 15 0
1 U
5697 0 0
2
45439.4 33
0
5 7415~
219 363 1497 0 4 22
0 144 143 142 141
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U20B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 15 0
1 U
3805 0 0
2
45439.4 34
0
8 2-In OR~
219 524 1528 0 3 22
0 146 145 90
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
5219 0 0
2
45439.4 35
0
8 2-In OR~
219 433 1646 0 3 22
0 135 134 145
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U23A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
3795 0 0
2
45439.4 36
0
8 3-In OR~
219 423 1506 0 4 22
0 141 139 136 146
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U22A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 17 0
1 U
3637 0 0
2
45439.4 37
0
8 4-In OR~
219 533 1320 0 5 22
0 111 103 110 101 91
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
3226 0 0
2
45439.4 38
0
9 Inverter~
13 198 1229 0 2 22
0 104 148
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
6966 0 0
2
45439.4 39
0
9 Inverter~
13 160 1211 0 2 22
0 101 149
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
9796 0 0
2
45439.4 40
0
9 2-In AND~
219 384 1220 0 3 22
0 149 148 147
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
5952 0 0
2
45439.4 41
0
9 2-In AND~
219 311 1194 0 3 22
0 104 101 150
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
3649 0 0
2
45439.4 42
0
9 Inverter~
13 97 1170 0 2 22
0 103 151
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
3716 0 0
2
45439.4 43
0
8 4-In OR~
219 568 1174 0 5 22
0 111 151 150 147 99
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
4797 0 0
2
45439.4 44
0
8 4-In OR~
219 575 1078 0 5 22
0 112 113 104 111 100
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U15A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
4681 0 0
2
5.90125e-315 5.32571e-315
0
6 74136~
219 127 769 0 3 22
0 104 101 152
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
9730 0 0
2
5.90125e-315 5.3568e-315
0
6 74136~
219 129 719 0 3 22
0 103 104 153
0
0 0 624 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9874 0 0
2
5.90125e-315 5.36716e-315
0
6 74136~
219 127 667 0 3 22
0 111 103 154
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
364 0 0
2
5.90125e-315 5.37752e-315
0
6 74136~
219 126 612 0 3 22
0 36 111 158
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3656 0 0
2
5.90125e-315 5.38788e-315
0
6 74136~
219 133 564 0 3 22
0 4 36 159
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3131 0 0
2
5.90125e-315 5.39306e-315
0
6 74136~
219 126 513 0 3 22
0 3 4 160
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6772 0 0
2
5.90125e-315 5.39824e-315
0
6 74136~
219 200 448 0 3 22
0 5 3 161
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9557 0 0
2
5.90125e-315 5.40342e-315
0
14 Logic Display~
6 1417 34 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5789 0 0
2
45439.4 45
0
14 Logic Display~
6 1382 24 0 1 2
10 92
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7328 0 0
2
45439.4 46
0
14 Logic Display~
6 1354 23 0 1 2
10 93
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4799 0 0
2
45439.4 47
0
14 Logic Display~
6 1332 23 0 1 2
10 94
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9196 0 0
2
45439.4 48
0
14 Logic Display~
6 1298 27 0 1 2
10 95
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3857 0 0
2
45439.4 49
0
14 Logic Display~
6 1273 31 0 1 2
10 96
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7125 0 0
2
45439.4 50
0
14 Logic Display~
6 1250 33 0 1 2
10 97
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
45439.4 51
0
14 Logic Display~
6 1215 34 0 1 2
10 98
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9821 0 0
2
45439.4 52
0
6 74136~
219 385 355 0 3 22
0 156 101 155
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3187 0 0
2
45439.4 53
0
6 74136~
219 335 331 0 3 22
0 157 104 156
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
762 0 0
2
45439.4 54
0
6 74136~
219 284 295 0 3 22
0 162 103 157
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
39 0 0
2
45439.4 55
0
6 74136~
219 237 266 0 3 22
0 163 111 162
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9450 0 0
2
45439.4 56
0
6 74136~
219 186 225 0 3 22
0 164 36 163
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3236 0 0
2
45439.4 57
0
7 74LS251
144 1023 801 0 14 29
0 214 215 216 217 218 155 28 152 6
7 8 17 219 16
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3321 0 0
2
5.90125e-315 5.4086e-315
0
7 74LS251
144 1027 699 0 14 29
0 220 221 222 223 224 156 84 153 6
7 8 17 225 92
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8879 0 0
2
5.90125e-315 5.41378e-315
0
7 74LS251
144 1027 599 0 14 29
0 226 227 228 229 230 157 85 154 6
7 8 17 231 93
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5433 0 0
2
5.90125e-315 5.41896e-315
0
7 74LS251
144 1027 492 0 14 29
0 232 233 234 235 236 162 86 158 6
7 8 17 237 94
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3679 0 0
2
5.90125e-315 5.42414e-315
0
7 74LS251
144 1028 389 0 14 29
0 238 239 240 241 242 163 90 159 6
7 8 17 243 95
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
9342 0 0
2
5.90125e-315 5.42933e-315
0
7 74LS251
144 1034 287 0 14 29
0 244 245 246 247 248 164 91 160 6
7 8 17 249 96
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3623 0 0
2
5.90125e-315 5.43192e-315
0
7 74LS251
144 1033 187 0 14 29
0 250 251 252 253 254 165 99 161 6
7 8 17 255 97
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3722 0 0
2
5.90125e-315 5.43451e-315
0
8 Hex Key~
166 1115 33 0 11 12
0 8 7 6 256 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8993 0 0
2
5.90125e-315 5.4371e-315
0
7 74LS251
144 1033 94 0 14 29
0 257 258 259 260 261 5 100 5 6
7 8 17 262 98
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-42 -37 -28 -29
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3723 0 0
2
5.90125e-315 5.43969e-315
0
8 Hex Key~
166 15 40 0 11 12
0 36 4 3 5 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6244 0 0
2
5.90125e-315 5.44487e-315
0
6 74136~
219 89 163 0 3 22
0 3 5 165
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-10 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6421 0 0
2
5.90125e-315 5.44746e-315
0
6 74136~
219 138 193 0 3 22
0 165 4 164
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7743 0 0
2
5.90125e-315 5.45264e-315
0
8 Hex Key~
166 52 42 0 11 12
0 101 104 103 111 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9840 0 0
2
5.90125e-315 5.45523e-315
0
362
0 1 3 0 0 4096 0 0 73 157 0 2
12 2411
243 2411
2 0 4 0 0 4096 0 74 0 0 156 2
539 2393
18 2393
1 0 5 0 0 4096 0 74 0 0 158 2
539 2384
6 2384
9 0 6 0 0 4096 0 6 0 0 40 2
1068 1223
1112 1223
0 10 7 0 0 4096 0 0 6 41 0 2
1118 1232
1068 1232
11 0 8 0 0 4096 0 6 0 0 42 2
1068 1241
1124 1241
1 0 5 0 0 4096 0 22 0 0 158 2
768 3281
6 3281
1 8 9 0 0 4224 0 1 3 0 0 3
1718 151
1561 151
1561 122
1 8 9 0 0 0 0 1 79 0 0 3
1718 151
1674 151
1674 127
1 9 2 0 0 8192 0 78 3 0 0 4
1596 20
1596 36
1540 36
1540 44
14 7 10 0 0 8320 0 4 3 0 0 3
1074 1489
1555 1489
1555 122
14 6 11 0 0 8320 0 5 3 0 0 3
1071 1391
1549 1391
1549 122
14 5 12 0 0 8320 0 6 3 0 0 3
1068 1286
1543 1286
1543 122
14 4 13 0 0 8320 0 7 3 0 0 3
1065 1176
1537 1176
1537 122
14 3 14 0 0 8320 0 8 3 0 0 3
1064 1061
1531 1061
1531 122
14 2 15 0 0 8320 0 9 3 0 0 3
1058 957
1525 957
1525 122
14 1 16 0 0 8192 0 155 3 0 0 3
1055 837
1519 837
1519 122
10 0 7 0 0 4096 0 8 0 0 41 2
1064 1007
1118 1007
11 0 8 0 0 4096 0 9 0 0 42 2
1058 912
1124 912
9 0 6 0 0 4096 0 8 0 0 40 2
1064 998
1112 998
11 0 8 0 0 0 0 8 0 0 42 2
1064 1016
1124 1016
9 0 6 0 0 4096 0 9 0 0 40 2
1058 894
1112 894
0 10 7 0 0 4096 0 0 9 41 0 2
1118 903
1058 903
12 0 17 0 0 4096 0 9 0 0 33 4
1064 921
1155 921
1155 922
1160 922
12 0 17 0 0 0 0 8 0 0 33 2
1070 1025
1160 1025
9 0 6 0 0 0 0 7 0 0 40 2
1065 1113
1112 1113
0 10 7 0 0 0 0 0 7 41 0 2
1118 1122
1065 1122
0 11 8 0 0 0 0 0 7 42 0 2
1124 1131
1065 1131
12 0 17 0 0 0 0 7 0 0 33 2
1071 1140
1160 1140
12 0 17 0 0 0 0 6 0 0 33 2
1074 1250
1160 1250
12 0 17 0 0 0 0 5 0 0 33 2
1077 1355
1160 1355
12 0 17 0 0 0 0 4 0 0 33 2
1080 1453
1160 1453
1 0 17 0 0 4224 0 2 0 0 0 2
1160 34
1160 1472
0 9 6 0 0 0 0 0 5 40 0 2
1112 1328
1071 1328
0 10 7 0 0 0 0 0 5 41 0 2
1118 1337
1071 1337
0 11 8 0 0 0 0 0 5 42 0 2
1124 1346
1071 1346
0 9 6 0 0 0 0 0 4 40 0 2
1112 1426
1074 1426
0 10 7 0 0 0 0 0 4 41 0 2
1118 1435
1074 1435
0 11 8 0 0 0 0 0 4 42 0 2
1124 1444
1074 1444
0 3 6 0 0 12416 0 0 162 0 0 4
1111 1456
1111 1426
1112 1426
1112 57
0 2 7 0 0 12416 0 0 162 0 0 4
1117 1456
1117 1435
1118 1435
1118 57
1 0 8 0 0 4224 0 162 0 0 0 4
1124 57
1124 1444
1123 1444
1123 1456
7 2 18 0 0 8320 0 4 11 0 0 3
1010 1480
984 1480
984 1893
7 2 19 0 0 8320 0 5 10 0 0 3
1007 1382
950 1382
950 1865
2 7 20 0 0 4224 0 38 6 0 0 3
924 1833
924 1277
1004 1277
2 1 21 0 0 4224 0 57 12 0 0 2
900 1796
900 1364
2 1 22 0 0 4224 0 60 13 0 0 2
881 1757
881 1240
1 2 23 0 0 4224 0 14 67 0 0 2
856 1236
856 1744
2 1 24 0 0 4224 0 68 15 0 0 2
824 1750
824 1238
7 2 25 0 0 8320 0 7 12 0 0 3
1001 1167
900 1167
900 1334
7 2 26 0 0 8320 0 8 13 0 0 3
1000 1052
881 1052
881 1210
7 2 27 0 0 8320 0 9 14 0 0 3
994 948
856 948
856 1206
7 2 28 0 0 8320 0 155 15 0 0 3
991 828
824 828
824 1208
5 1 29 0 0 8320 0 22 11 0 0 3
818 3294
984 3294
984 1923
1 5 30 0 0 4224 0 10 30 0 0 3
950 1895
950 3134
749 3134
3 3 31 0 0 4224 0 22 20 0 0 4
768 3299
447 3299
447 3354
439 3354
3 4 32 0 0 4224 0 19 22 0 0 4
538 3394
760 3394
760 3308
768 3308
3 2 33 0 0 12416 0 21 22 0 0 4
366 3307
394 3307
394 3290
768 3290
1 0 4 0 0 0 0 16 0 0 156 2
249 3403
18 3403
1 0 3 0 0 0 0 17 0 0 157 2
135 3345
12 3345
2 2 34 0 0 4224 0 16 19 0 0 2
285 3403
493 3403
2 1 35 0 0 4224 0 17 20 0 0 2
171 3345
394 3345
1 0 3 0 0 4096 0 19 0 0 157 2
493 3385
12 3385
2 0 4 0 0 0 0 20 0 0 156 2
394 3363
18 3363
1 0 36 0 0 4096 0 18 0 0 155 4
185 3316
29 3316
29 3317
24 3317
2 2 37 0 0 4224 0 18 21 0 0 2
221 3316
321 3316
1 0 4 0 0 0 0 21 0 0 156 2
321 3298
18 3298
1 0 4 0 0 0 0 23 0 0 156 2
169 3253
18 3253
2 2 38 0 0 4224 0 23 27 0 0 2
205 3253
442 3253
1 0 3 0 0 0 0 27 0 0 157 2
442 3235
12 3235
1 0 36 0 0 4096 0 24 0 0 155 2
217 3207
24 3207
2 2 39 0 0 4224 0 24 28 0 0 2
253 3207
400 3207
1 0 3 0 0 0 0 28 0 0 157 2
400 3189
12 3189
1 0 36 0 0 4096 0 25 0 0 155 2
220 3162
24 3162
1 0 4 0 0 0 0 26 0 0 156 2
182 3144
18 3144
2 2 40 0 0 4224 0 29 25 0 0 2
366 3162
256 3162
2 1 41 0 0 4224 0 26 29 0 0 2
218 3144
366 3144
3 4 42 0 0 12416 0 27 30 0 0 4
487 3244
578 3244
578 3148
699 3148
3 3 43 0 0 12416 0 28 30 0 0 4
445 3198
514 3198
514 3139
699 3139
3 2 44 0 0 8320 0 29 30 0 0 3
411 3153
411 3130
699 3130
1 0 5 0 0 0 0 30 0 0 158 2
699 3121
6 3121
1 0 36 0 0 0 0 31 0 0 155 4
133 3090
29 3090
29 3091
24 3091
1 0 4 0 0 0 0 35 0 0 156 2
357 3072
18 3072
2 2 45 0 0 4224 0 31 35 0 0 2
169 3090
357 3090
1 0 36 0 0 0 0 32 0 0 155 4
115 3040
29 3040
29 3041
24 3041
1 0 4 0 0 0 0 33 0 0 156 2
201 3031
18 3031
1 0 3 0 0 0 0 34 0 0 157 2
282 3022
12 3022
3 2 46 0 0 4224 0 36 32 0 0 2
356 3040
151 3040
2 2 47 0 0 4224 0 36 33 0 0 2
356 3031
237 3031
2 1 48 0 0 4224 0 34 36 0 0 2
318 3022
356 3022
2 3 49 0 0 12416 0 37 35 0 0 4
714 3062
567 3062
567 3081
402 3081
4 1 50 0 0 4224 0 36 37 0 0 4
401 3031
706 3031
706 3044
714 3044
3 1 51 0 0 8320 0 37 38 0 0 3
760 3053
924 3053
924 1863
1 0 36 0 0 0 0 39 0 0 155 4
125 2967
29 2967
29 2968
24 2968
1 0 5 0 0 0 0 40 0 0 158 2
222 2949
6 2949
2 1 52 0 0 4224 0 40 50 0 0 2
258 2949
359 2949
3 2 53 0 0 4224 0 50 39 0 0 2
359 2967
161 2967
2 0 4 0 0 0 0 50 0 0 156 2
359 2958
18 2958
1 0 5 0 0 0 0 42 0 0 158 2
199 2900
6 2900
1 0 3 0 0 0 0 41 0 0 157 2
139 2909
12 2909
3 0 4 0 0 0 0 51 0 0 156 2
358 2918
18 2918
2 2 54 0 0 4224 0 51 41 0 0 2
358 2909
175 2909
2 1 55 0 0 4224 0 42 51 0 0 2
235 2900
358 2900
1 0 4 0 0 0 0 43 0 0 156 2
252 2865
18 2865
1 0 3 0 0 0 0 44 0 0 157 2
178 2856
12 2856
2 2 56 0 0 4224 0 52 44 0 0 2
357 2856
214 2856
2 3 57 0 0 4224 0 43 52 0 0 2
288 2865
357 2865
1 0 5 0 0 0 0 52 0 0 158 2
357 2847
6 2847
1 0 4 0 0 0 0 45 0 0 156 2
132 2804
18 2804
2 2 58 0 0 4224 0 45 53 0 0 2
168 2804
295 2804
3 0 36 0 0 4096 0 53 0 0 155 2
295 2813
24 2813
1 0 3 0 0 0 0 53 0 0 157 2
295 2795
12 2795
1 3 59 0 0 4224 0 49 56 0 0 4
716 2834
628 2834
628 2786
606 2786
4 2 60 0 0 12416 0 55 49 0 0 4
610 2884
625 2884
625 2852
716 2852
3 4 61 0 0 12416 0 55 50 0 0 4
564 2893
490 2893
490 2958
404 2958
4 2 62 0 0 12416 0 51 55 0 0 4
403 2909
440 2909
440 2884
565 2884
1 4 63 0 0 4224 0 55 52 0 0 4
564 2875
410 2875
410 2856
402 2856
2 4 64 0 0 4224 0 56 53 0 0 4
560 2795
410 2795
410 2804
340 2804
4 1 65 0 0 4224 0 54 56 0 0 4
338 2753
552 2753
552 2777
560 2777
2 3 66 0 0 4224 0 46 54 0 0 2
206 2762
293 2762
2 2 67 0 0 4224 0 54 47 0 0 2
293 2753
76 2753
2 1 68 0 0 4224 0 48 54 0 0 2
118 2744
293 2744
1 0 36 0 0 0 0 46 0 0 155 2
170 2762
24 2762
1 0 4 0 0 0 0 47 0 0 156 2
40 2753
18 2753
1 0 3 0 0 0 0 48 0 0 157 2
82 2744
12 2744
3 1 69 0 0 8320 0 49 57 0 0 3
762 2843
900 2843
900 1826
5 1 70 0 0 8320 0 59 60 0 0 3
607 2684
881 2684
881 1787
1 0 4 0 0 0 0 58 0 0 156 2
197 2689
18 2689
2 3 71 0 0 4224 0 58 59 0 0 2
233 2689
557 2689
4 0 36 0 0 4096 0 59 0 0 155 2
557 2698
24 2698
2 0 3 0 0 4096 0 59 0 0 157 2
557 2680
12 2680
1 0 5 0 0 0 0 59 0 0 158 2
557 2671
6 2671
1 5 72 0 0 4224 0 67 66 0 0 3
856 1774
856 2554
594 2554
1 0 36 0 0 0 0 61 0 0 155 2
112 2628
24 2628
1 0 4 0 0 0 0 62 0 0 156 2
160 2610
18 2610
4 3 73 0 0 12416 0 66 63 0 0 4
544 2568
480 2568
480 2619
307 2619
3 3 74 0 0 12416 0 64 66 0 0 4
370 2573
446 2573
446 2559
544 2559
2 2 75 0 0 4224 0 61 63 0 0 2
148 2628
262 2628
1 2 76 0 0 4224 0 63 62 0 0 2
262 2610
196 2610
0 2 36 0 0 0 0 0 64 155 0 2
24 2582
325 2582
1 0 4 0 0 0 0 64 0 0 156 2
325 2564
18 2564
2 2 77 0 0 4224 0 65 66 0 0 2
156 2550
544 2550
1 0 3 0 0 0 0 65 0 0 157 2
120 2550
12 2550
1 0 5 0 0 0 0 66 0 0 158 2
544 2541
6 2541
5 1 78 0 0 8320 0 74 68 0 0 3
589 2397
824 2397
824 1780
4 4 79 0 0 4224 0 72 74 0 0 4
382 2461
480 2461
480 2411
539 2411
1 0 36 0 0 0 0 69 0 0 155 2
174 2470
24 2470
1 0 4 0 0 0 0 70 0 0 156 2
90 2461
18 2461
1 0 3 0 0 0 0 71 0 0 157 2
139 2452
12 2452
2 1 80 0 0 4224 0 71 72 0 0 2
175 2452
337 2452
2 2 81 0 0 4224 0 72 70 0 0 2
337 2461
126 2461
2 3 82 0 0 4224 0 69 72 0 0 2
210 2470
337 2470
2 0 36 0 0 0 0 73 0 0 155 2
243 2429
24 2429
3 3 83 0 0 12416 0 73 74 0 0 4
288 2420
389 2420
389 2402
539 2402
0 1 36 0 0 4224 0 0 164 0 0 2
24 3413
24 64
2 0 4 0 0 4224 0 164 0 0 0 2
18 64
18 3413
0 3 3 0 0 4224 0 0 164 0 0 2
12 3413
12 64
4 0 5 0 0 4224 0 164 0 0 0 2
6 64
6 3413
2 7 84 0 0 4224 0 75 156 0 0 3
787 1207
787 726
995 726
7 2 85 0 0 8320 0 157 76 0 0 3
995 626
758 626
758 1205
2 7 86 0 0 4224 0 77 158 0 0 3
726 1202
726 519
995 519
1 5 87 0 0 4224 0 75 99 0 0 3
787 1237
787 2173
595 2173
5 1 88 0 0 8320 0 107 76 0 0 3
587 1976
758 1976
758 1235
1 3 89 0 0 4224 0 77 86 0 0 3
726 1232
726 1759
566 1759
7 3 90 0 0 8320 0 159 124 0 0 4
996 416
710 416
710 1528
557 1528
7 5 91 0 0 8320 0 160 127 0 0 6
1002 314
696 314
696 1319
574 1319
574 1320
566 1320
14 7 92 0 0 4096 0 156 79 0 0 3
1059 735
1668 735
1668 127
6 14 93 0 0 8320 0 79 157 0 0 3
1662 127
1662 635
1059 635
14 5 94 0 0 4224 0 158 79 0 0 3
1059 528
1656 528
1656 127
4 14 95 0 0 8320 0 79 159 0 0 3
1650 127
1650 425
1060 425
14 3 96 0 0 4224 0 160 79 0 0 3
1066 323
1644 323
1644 127
2 14 97 0 0 8320 0 79 161 0 0 3
1638 127
1638 223
1065 223
14 1 98 0 0 4224 0 163 79 0 0 3
1065 130
1632 130
1632 127
5 7 99 0 0 8320 0 133 161 0 0 4
601 1174
682 1174
682 214
1001 214
5 7 100 0 0 8320 0 134 163 0 0 4
608 1078
664 1078
664 121
1001 121
9 1 2 0 0 8320 0 79 78 0 0 4
1653 49
1653 35
1596 35
1596 20
1 0 101 0 0 4096 0 80 0 0 255 2
114 1840
61 1840
2 2 102 0 0 4224 0 80 84 0 0 2
150 1840
191 1840
1 0 103 0 0 4096 0 81 0 0 257 2
195 1741
49 1741
1 0 104 0 0 4096 0 82 0 0 256 2
142 1750
55 1750
2 1 105 0 0 4224 0 81 85 0 0 2
231 1741
249 1741
2 2 106 0 0 4224 0 82 85 0 0 2
178 1750
249 1750
1 0 101 0 0 0 0 83 0 0 255 2
95 1759
61 1759
2 3 107 0 0 4224 0 83 85 0 0 2
131 1759
249 1759
4 1 108 0 0 4224 0 85 86 0 0 2
294 1750
520 1750
3 2 109 0 0 4224 0 84 86 0 0 4
236 1831
398 1831
398 1768
520 1768
1 0 104 0 0 4096 0 84 0 0 256 2
191 1822
55 1822
4 0 101 0 0 4096 0 127 0 0 255 2
516 1334
61 1334
1 0 104 0 0 0 0 87 0 0 256 2
188 1325
55 1325
2 3 110 0 0 4224 0 87 127 0 0 2
224 1325
516 1325
2 0 103 0 0 4096 0 127 0 0 257 2
516 1316
49 1316
1 0 111 0 0 4096 0 127 0 0 258 2
516 1307
43 1307
1 0 101 0 0 0 0 88 0 0 255 2
302 938
61 938
2 0 103 0 0 0 0 88 0 0 257 2
302 956
49 956
3 1 112 0 0 12416 0 88 134 0 0 4
347 947
433 947
433 1065
558 1065
4 0 111 0 0 4096 0 134 0 0 258 2
558 1092
43 1092
3 0 104 0 0 4096 0 134 0 0 256 2
558 1083
55 1083
2 4 113 0 0 4224 0 134 92 0 0 4
558 1074
378 1074
378 1000
370 1000
1 0 101 0 0 0 0 89 0 0 255 2
105 1009
61 1009
1 0 104 0 0 0 0 90 0 0 256 2
148 1000
55 1000
1 0 103 0 0 0 0 91 0 0 257 2
188 991
49 991
3 2 114 0 0 4224 0 92 89 0 0 2
325 1009
141 1009
2 2 115 0 0 4224 0 92 90 0 0 2
325 1000
184 1000
2 1 116 0 0 4224 0 91 92 0 0 2
224 991
325 991
1 0 103 0 0 0 0 96 0 0 257 2
378 2250
49 2250
1 0 104 0 0 0 0 93 0 0 256 2
200 2268
55 2268
2 2 117 0 0 4224 0 93 96 0 0 2
236 2268
378 2268
2 0 104 0 0 0 0 97 0 0 256 2
321 2233
55 2233
1 0 103 0 0 0 0 94 0 0 257 2
191 2215
49 2215
2 1 118 0 0 4224 0 94 97 0 0 2
227 2215
321 2215
2 0 104 0 0 0 0 98 0 0 256 2
370 2190
55 2190
1 0 101 0 0 0 0 95 0 0 255 2
205 2172
61 2172
2 1 119 0 0 4224 0 95 98 0 0 2
241 2172
370 2172
4 3 120 0 0 12416 0 99 96 0 0 4
545 2187
516 2187
516 2259
423 2259
3 3 121 0 0 12416 0 99 97 0 0 4
545 2178
470 2178
470 2224
366 2224
3 2 122 0 0 12416 0 98 99 0 0 4
415 2181
451 2181
451 2169
545 2169
1 0 111 0 0 0 0 99 0 0 258 2
545 2160
43 2160
3 4 123 0 0 4224 0 104 107 0 0 4
392 2070
529 2070
529 1990
537 1990
3 3 124 0 0 12416 0 105 107 0 0 4
388 2018
421 2018
421 1981
537 1981
1 0 104 0 0 0 0 100 0 0 256 2
218 2079
55 2079
1 0 103 0 0 0 0 105 0 0 257 2
343 2009
49 2009
2 2 125 0 0 4224 0 100 104 0 0 2
254 2079
347 2079
1 0 103 0 0 0 0 104 0 0 257 2
347 2061
49 2061
1 0 101 0 0 0 0 101 0 0 255 2
218 2027
61 2027
2 2 126 0 0 4224 0 101 105 0 0 2
254 2027
343 2027
3 2 127 0 0 12416 0 106 107 0 0 4
330 1982
381 1982
381 1972
537 1972
2 2 128 0 0 4224 0 106 103 0 0 2
285 1991
165 1991
2 1 129 0 0 4224 0 102 106 0 0 2
222 1973
285 1973
1 0 101 0 0 0 0 103 0 0 255 2
129 1991
61 1991
1 0 104 0 0 0 0 102 0 0 256 2
186 1973
55 1973
1 0 111 0 0 0 0 107 0 0 258 2
537 1963
43 1963
1 0 101 0 0 0 0 108 0 0 255 2
127 1685
61 1685
2 3 130 0 0 4224 0 108 119 0 0 2
163 1685
341 1685
2 0 104 0 0 0 0 119 0 0 256 2
341 1676
55 1676
1 0 111 0 0 0 0 109 0 0 258 2
183 1667
43 1667
2 1 131 0 0 4224 0 109 119 0 0 2
219 1667
341 1667
1 0 103 0 0 0 0 110 0 0 257 2
152 1622
49 1622
2 2 132 0 0 4224 0 110 122 0 0 2
188 1622
299 1622
1 0 111 0 0 0 0 111 0 0 258 2
75 1613
43 1613
2 1 133 0 0 4224 0 111 122 0 0 2
111 1613
299 1613
3 0 104 0 0 0 0 122 0 0 256 2
299 1631
55 1631
4 2 134 0 0 4224 0 119 125 0 0 4
386 1676
412 1676
412 1655
420 1655
4 1 135 0 0 4224 0 122 125 0 0 4
344 1622
412 1622
412 1637
420 1637
4 3 136 0 0 8320 0 120 126 0 0 4
387 1568
402 1568
402 1515
410 1515
1 0 104 0 0 0 0 112 0 0 256 2
235 1577
55 1577
1 0 103 0 0 0 0 113 0 0 257 2
156 1568
49 1568
2 3 137 0 0 4224 0 112 120 0 0 2
271 1577
342 1577
2 2 138 0 0 4224 0 113 120 0 0 2
192 1568
342 1568
1 0 111 0 0 0 0 120 0 0 258 2
342 1559
43 1559
3 0 101 0 0 0 0 121 0 0 255 2
299 1543
61 1543
1 0 104 0 0 0 0 114 0 0 256 2
206 1534
55 1534
4 2 139 0 0 4224 0 121 126 0 0 4
344 1534
381 1534
381 1506
411 1506
2 2 140 0 0 4224 0 114 121 0 0 2
242 1534
299 1534
0 1 103 0 0 0 0 0 121 257 0 2
49 1525
299 1525
1 4 101 0 0 4224 0 167 115 0 0 4
61 66
61 1840
62 1840
62 2280
2 3 104 0 0 4224 0 167 115 0 0 4
55 66
55 1822
56 1822
56 2280
3 2 103 0 0 4224 0 167 115 0 0 4
49 66
49 1741
50 1741
50 2280
4 1 111 0 0 4224 0 167 115 0 0 4
43 66
43 1307
44 1307
44 2280
4 1 141 0 0 4224 0 123 126 0 0 2
384 1497
410 1497
2 3 142 0 0 4224 0 116 123 0 0 2
203 1506
339 1506
2 2 143 0 0 4224 0 123 117 0 0 2
339 1497
252 1497
2 1 144 0 0 4224 0 118 123 0 0 2
299 1488
339 1488
1 1 101 0 0 0 0 167 116 0 0 3
61 66
61 1506
167 1506
2 1 104 0 0 0 0 167 117 0 0 3
55 66
55 1497
216 1497
3 1 103 0 0 0 0 167 118 0 0 3
49 66
49 1488
263 1488
2 3 145 0 0 8320 0 124 125 0 0 4
511 1537
490 1537
490 1646
466 1646
4 1 146 0 0 4224 0 126 124 0 0 4
456 1506
489 1506
489 1519
511 1519
3 4 147 0 0 12416 0 130 133 0 0 4
405 1220
471 1220
471 1188
551 1188
2 2 148 0 0 4224 0 130 128 0 0 2
360 1229
219 1229
2 1 149 0 0 4224 0 129 130 0 0 2
181 1211
360 1211
2 1 104 0 0 0 0 167 128 0 0 3
55 66
55 1229
183 1229
1 1 101 0 0 0 0 167 129 0 0 3
61 66
61 1211
145 1211
3 3 150 0 0 12416 0 131 133 0 0 4
332 1194
368 1194
368 1179
551 1179
1 2 101 0 0 0 0 167 131 0 0 3
61 66
61 1203
287 1203
2 1 104 0 0 0 0 167 131 0 0 3
55 66
55 1185
287 1185
2 2 151 0 0 4224 0 132 133 0 0 2
118 1170
551 1170
3 1 103 0 0 0 0 167 132 0 0 3
49 66
49 1170
82 1170
4 1 111 0 0 0 0 167 133 0 0 3
43 66
43 1161
551 1161
4 1 5 0 0 0 0 164 141 0 0 3
6 64
6 439
184 439
3 8 152 0 0 4224 0 135 155 0 0 4
160 769
603 769
603 837
991 837
3 8 153 0 0 16512 0 136 156 0 0 5
162 719
162 724
577 724
577 735
995 735
3 8 154 0 0 12416 0 137 157 0 0 4
160 667
566 667
566 635
995 635
3 6 155 0 0 8320 0 150 155 0 0 4
418 355
528 355
528 819
991 819
3 6 156 0 0 12416 0 151 156 0 0 4
368 331
537 331
537 717
995 717
3 6 157 0 0 12416 0 152 157 0 0 4
317 295
550 295
550 617
995 617
1 2 101 0 0 0 0 167 135 0 0 3
61 66
61 778
111 778
2 1 104 0 0 0 0 167 135 0 0 3
55 66
55 760
111 760
2 2 104 0 0 0 0 136 167 0 0 3
113 728
55 728
55 66
3 1 103 0 0 0 0 167 136 0 0 3
49 66
49 710
113 710
3 2 103 0 0 0 0 167 137 0 0 3
49 66
49 676
111 676
4 1 111 0 0 0 0 167 137 0 0 3
43 66
43 658
111 658
3 8 158 0 0 4224 0 138 158 0 0 4
159 612
605 612
605 528
995 528
4 2 111 0 0 0 0 167 138 0 0 3
43 66
43 621
110 621
1 1 36 0 0 0 0 164 138 0 0 3
24 64
24 603
110 603
3 8 159 0 0 4224 0 139 159 0 0 4
166 564
599 564
599 425
996 425
3 8 160 0 0 4224 0 140 160 0 0 4
159 513
592 513
592 323
1002 323
3 8 161 0 0 12416 0 141 161 0 0 4
233 448
583 448
583 223
1001 223
2 1 36 0 0 0 0 139 164 0 0 3
117 573
24 573
24 64
2 1 4 0 0 0 0 164 139 0 0 3
18 64
18 555
117 555
2 2 4 0 0 0 0 140 164 0 0 3
110 522
18 522
18 64
3 1 3 0 0 0 0 164 140 0 0 3
12 64
12 504
110 504
2 3 3 0 0 0 0 141 164 0 0 3
184 457
12 457
12 64
3 6 162 0 0 12416 0 153 158 0 0 4
270 266
518 266
518 510
995 510
3 6 163 0 0 12416 0 154 159 0 0 4
219 225
501 225
501 407
996 407
3 6 164 0 0 12416 0 166 160 0 0 4
171 193
511 193
511 305
1002 305
3 6 165 0 0 12416 0 165 161 0 0 4
122 163
516 163
516 205
1001 205
4 8 5 0 0 0 0 164 163 0 0 3
6 64
6 130
1001 130
4 6 5 0 0 0 0 164 163 0 0 3
6 64
6 112
1001 112
14 1 16 0 0 8320 0 155 142 0 0 3
1055 837
1417 837
1417 52
14 1 92 0 0 8320 0 156 143 0 0 3
1059 735
1382 735
1382 42
14 1 93 0 0 0 0 157 144 0 0 3
1059 635
1354 635
1354 41
14 1 94 0 0 0 0 158 145 0 0 3
1059 528
1332 528
1332 41
14 1 95 0 0 0 0 159 146 0 0 3
1060 425
1298 425
1298 45
14 1 96 0 0 0 0 160 147 0 0 3
1066 323
1273 323
1273 49
14 1 97 0 0 0 0 161 148 0 0 3
1065 223
1250 223
1250 51
14 1 98 0 0 0 0 163 149 0 0 3
1065 130
1215 130
1215 52
2 1 101 0 0 0 0 150 167 0 0 3
369 364
61 364
61 66
3 1 156 0 0 0 0 151 150 0 0 4
368 331
366 331
366 346
369 346
2 2 104 0 0 0 0 151 167 0 0 3
319 340
55 340
55 66
3 1 157 0 0 0 0 152 151 0 0 3
317 295
317 322
319 322
2 3 103 0 0 0 0 152 167 0 0 3
268 304
49 304
49 66
3 1 162 0 0 0 0 153 152 0 0 3
270 266
268 266
268 286
4 2 111 0 0 0 0 167 153 0 0 3
43 66
43 275
221 275
3 1 163 0 0 0 0 154 153 0 0 4
219 225
220 225
220 257
221 257
1 2 36 0 0 0 0 164 154 0 0 3
24 64
24 234
170 234
3 1 164 0 0 0 0 166 154 0 0 4
171 193
169 193
169 216
170 216
2 2 4 0 0 0 0 164 166 0 0 3
18 64
18 202
122 202
12 1 17 0 0 0 0 155 2 0 0 3
1061 801
1160 801
1160 34
12 1 17 0 0 0 0 156 2 0 0 3
1065 699
1160 699
1160 34
12 1 17 0 0 0 0 157 2 0 0 3
1065 599
1160 599
1160 34
12 1 17 0 0 0 0 158 2 0 0 3
1065 492
1160 492
1160 34
12 1 17 0 0 0 0 159 2 0 0 3
1066 389
1160 389
1160 34
12 1 17 0 0 0 0 160 2 0 0 3
1072 287
1160 287
1160 34
12 1 17 0 0 0 0 161 2 0 0 3
1071 187
1160 187
1160 34
1 12 17 0 0 0 0 2 163 0 0 3
1160 34
1160 94
1071 94
9 3 6 0 0 0 0 157 162 0 0 3
1059 572
1112 572
1112 57
9 3 6 0 0 0 0 156 162 0 0 3
1059 672
1112 672
1112 57
3 9 6 0 0 0 0 162 155 0 0 3
1112 57
1112 774
1055 774
10 2 7 0 0 0 0 155 162 0 0 3
1055 783
1118 783
1118 57
10 2 7 0 0 0 0 156 162 0 0 3
1059 681
1118 681
1118 57
2 10 7 0 0 0 0 162 157 0 0 3
1118 57
1118 581
1059 581
11 1 8 0 0 0 0 155 162 0 0 3
1055 792
1124 792
1124 57
11 1 8 0 0 0 0 156 162 0 0 3
1059 690
1124 690
1124 57
11 1 8 0 0 0 0 157 162 0 0 3
1059 590
1124 590
1124 57
9 3 6 0 0 0 0 158 162 0 0 3
1059 465
1112 465
1112 57
9 3 6 0 0 0 0 159 162 0 0 3
1060 362
1112 362
1112 57
2 10 7 0 0 0 0 162 158 0 0 3
1118 57
1118 474
1059 474
2 10 7 0 0 0 0 162 159 0 0 3
1118 57
1118 371
1060 371
11 1 8 0 0 0 0 158 162 0 0 3
1059 483
1124 483
1124 57
1 11 8 0 0 0 0 162 159 0 0 3
1124 57
1124 380
1060 380
1 11 8 0 0 0 0 162 160 0 0 3
1124 57
1124 278
1066 278
10 2 7 0 0 0 0 160 162 0 0 3
1066 269
1118 269
1118 57
3 9 6 0 0 0 0 162 160 0 0 3
1112 57
1112 260
1066 260
11 1 8 0 0 0 0 161 162 0 0 3
1065 178
1124 178
1124 57
2 10 7 0 0 0 0 162 161 0 0 3
1118 57
1118 169
1065 169
9 3 6 0 0 0 0 161 162 0 0 3
1065 160
1112 160
1112 57
3 9 6 0 0 0 0 162 163 0 0 3
1112 57
1112 67
1065 67
2 10 7 0 0 0 0 162 163 0 0 3
1118 57
1118 76
1065 76
1 11 8 0 0 0 0 162 163 0 0 3
1124 57
1124 85
1065 85
3 1 3 0 0 0 0 164 165 0 0 3
12 64
12 154
73 154
4 2 5 0 0 0 0 164 165 0 0 3
6 64
6 172
73 172
3 1 165 0 0 0 0 165 166 0 0 2
122 163
122 184
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
949 -8 1096 53
959 2 1085 47
52 0=Binario->Grey
1=Binario->Displey
2=Grey->Binario
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
