CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
370 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 1160 22 0 1 11
0 6
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
45434.7 0
0
7 74LS251
144 1030 946 0 14 29
0 30 31 32 33 34 35 36 14 11
12 13 6 37 5
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
6369 0 0
2
45434.7 0
0
7 74LS251
144 1027 830 0 14 29
0 38 39 40 41 42 43 44 15 11
12 13 6 45 4
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
45434.7 0
0
7 74LS251
144 1028 722 0 14 29
0 46 47 48 49 50 51 52 16 11
12 13 6 53 3
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
7100 0 0
2
45434.7 0
0
7 74LS251
144 1028 615 0 14 29
0 54 55 56 57 58 59 60 17 11
12 13 6 61 2
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3820 0 0
2
45434.7 0
0
7 74LS251
144 1028 389 0 14 29
0 62 63 64 65 66 67 68 18 11
12 13 6 69 7
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
7678 0 0
2
45434.7 0
0
7 74LS251
144 1034 287 0 14 29
0 70 71 72 73 74 75 76 19 11
12 13 6 77 8
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
961 0 0
2
45434.7 0
0
7 74LS251
144 1033 187 0 14 29
0 78 79 80 81 82 83 84 20 11
12 13 6 85 9
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3178 0 0
2
45434.7 0
0
8 Hex Key~
166 1115 33 0 11 12
0 13 12 11 86 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
3409 0 0
2
45434.6 0
0
7 74LS251
144 1033 94 0 14 29
0 87 88 89 90 91 92 93 21 11
12 13 6 94 10
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3951 0 0
2
45434.6 0
0
12 Hex Display~
7 1417 45 0 16 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8885 0 0
2
45434.6 0
0
6 74136~
219 447 377 0 3 22
0 15 22 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3780 0 0
2
45434.6 0
0
6 74136~
219 400 347 0 3 22
0 16 23 15
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9265 0 0
2
45434.6 0
0
6 74136~
219 345 312 0 3 22
0 17 24 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9442 0 0
2
45434.6 0
0
6 74136~
219 301 286 0 3 22
0 26 25 17
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9424 0 0
2
45434.6 0
0
6 74136~
219 247 258 0 3 22
0 18 27 26
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9968 0 0
2
45434.6 0
0
6 74136~
219 190 230 0 3 22
0 19 28 18
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9281 0 0
2
45434.6 0
0
8 Hex Key~
166 16 44 0 11 12
0 27 28 29 21 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
8464 0 0
2
45434.6 0
0
6 74136~
219 89 163 0 3 22
0 29 21 20
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7168 0 0
2
45434.6 0
0
12 Hex Display~
7 1368 49 0 16 19
10 7 8 9 10 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3171 0 0
2
45434.6 0
0
6 74136~
219 138 194 0 3 22
0 20 29 19
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4139 0 0
2
45434.6 0
0
8 Hex Key~
166 52 42 0 11 12
0 22 23 24 25 0 0 0 0 0
8 56
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
6435 0 0
2
45434.6 0
0
68
14 4 2 0 0 8320 0 5 11 0 0 3
1060 651
1408 651
1408 69
14 3 3 0 0 8320 0 4 11 0 0 3
1060 758
1414 758
1414 69
14 2 4 0 0 8320 0 3 11 0 0 3
1059 866
1420 866
1420 69
14 1 5 0 0 8320 0 2 11 0 0 3
1062 982
1426 982
1426 69
12 1 6 0 0 8320 0 2 1 0 0 3
1068 946
1160 946
1160 34
12 1 6 0 0 0 0 3 1 0 0 3
1065 830
1160 830
1160 34
12 1 6 0 0 0 0 4 1 0 0 3
1066 722
1160 722
1160 34
12 1 6 0 0 0 0 5 1 0 0 3
1066 615
1160 615
1160 34
0 1 6 0 0 0 0 0 1 0 0 3
1067 505
1160 505
1160 34
12 1 6 0 0 0 0 6 1 0 0 3
1066 389
1160 389
1160 34
12 1 6 0 0 0 0 7 1 0 0 3
1072 287
1160 287
1160 34
12 1 6 0 0 0 0 8 1 0 0 3
1071 187
1160 187
1160 34
1 12 6 0 0 16 0 1 10 0 0 3
1160 34
1160 94
1071 94
14 1 7 0 0 8320 0 6 20 0 0 3
1060 425
1377 425
1377 73
14 2 8 0 0 4224 0 7 20 0 0 3
1066 323
1371 323
1371 73
14 3 9 0 0 4224 0 8 20 0 0 3
1065 223
1365 223
1365 73
14 4 10 0 0 4224 0 10 20 0 0 3
1065 130
1359 130
1359 73
9 3 11 0 0 8192 0 4 9 0 0 3
1060 695
1112 695
1112 57
9 3 11 0 0 8192 0 3 9 0 0 3
1059 803
1112 803
1112 57
3 9 11 0 0 4224 0 9 2 0 0 3
1112 57
1112 919
1062 919
10 2 12 0 0 8320 0 2 9 0 0 3
1062 928
1118 928
1118 57
10 2 12 0 0 0 0 3 9 0 0 3
1059 812
1118 812
1118 57
2 10 12 0 0 0 0 9 4 0 0 3
1118 57
1118 704
1060 704
11 1 13 0 0 8320 0 2 9 0 0 3
1062 937
1124 937
1124 57
11 1 13 0 0 0 0 3 9 0 0 3
1059 821
1124 821
1124 57
11 1 13 0 0 0 0 4 9 0 0 3
1060 713
1124 713
1124 57
9 3 11 0 0 0 0 5 9 0 0 3
1060 588
1112 588
1112 57
0 3 11 0 0 0 0 0 9 0 0 3
1061 478
1112 478
1112 57
9 3 11 0 0 0 0 6 9 0 0 3
1060 362
1112 362
1112 57
0 2 12 0 0 0 0 0 9 0 0 3
1061 487
1118 487
1118 57
2 10 12 0 0 0 0 9 5 0 0 3
1118 57
1118 597
1060 597
2 10 12 0 0 0 0 9 6 0 0 3
1118 57
1118 371
1060 371
11 1 13 0 0 0 0 5 9 0 0 3
1060 606
1124 606
1124 57
0 1 13 0 0 0 0 0 9 0 0 3
1061 496
1124 496
1124 57
1 11 13 0 0 0 0 9 6 0 0 3
1124 57
1124 380
1060 380
3 8 14 0 0 8320 0 12 2 0 0 4
480 377
759 377
759 982
998 982
3 8 15 0 0 8320 0 13 3 0 0 4
433 347
778 347
778 866
995 866
3 8 16 0 0 8320 0 14 4 0 0 4
378 312
796 312
796 758
996 758
3 8 17 0 0 4224 0 15 5 0 0 4
334 286
822 286
822 651
996 651
3 8 18 0 0 4224 0 17 6 0 0 4
223 230
861 230
861 425
996 425
3 8 19 0 0 4224 0 21 7 0 0 4
171 194
879 194
879 323
1002 323
3 8 20 0 0 4224 0 19 8 0 0 4
122 163
897 163
897 223
1001 223
4 8 21 0 0 8320 0 18 10 0 0 3
7 68
7 130
1001 130
1 11 13 0 0 0 0 9 7 0 0 3
1124 57
1124 278
1066 278
10 2 12 0 0 0 0 7 9 0 0 3
1066 269
1118 269
1118 57
3 9 11 0 0 0 0 9 7 0 0 3
1112 57
1112 260
1066 260
11 1 13 0 0 0 0 8 9 0 0 3
1065 178
1124 178
1124 57
2 10 12 0 0 0 0 9 8 0 0 3
1118 57
1118 169
1065 169
9 3 11 0 0 0 0 8 9 0 0 3
1065 160
1112 160
1112 57
3 9 11 0 0 0 0 9 10 0 0 3
1112 57
1112 67
1065 67
2 10 12 0 0 0 0 9 10 0 0 3
1118 57
1118 76
1065 76
1 11 13 0 0 0 0 9 10 0 0 3
1124 57
1124 85
1065 85
2 1 22 0 0 4224 0 12 22 0 0 3
431 386
61 386
61 66
3 1 15 0 0 0 0 13 12 0 0 3
433 347
433 368
431 368
2 2 23 0 0 8320 0 22 13 0 0 3
55 66
55 356
384 356
2 3 24 0 0 4224 0 14 22 0 0 3
329 321
49 321
49 66
3 1 16 0 0 0 0 14 13 0 0 4
378 312
388 312
388 338
384 338
3 1 17 0 0 0 0 15 14 0 0 4
334 286
332 286
332 303
329 303
4 2 25 0 0 8320 0 22 15 0 0 3
43 66
43 295
285 295
3 1 26 0 0 8320 0 16 15 0 0 4
280 258
281 258
281 277
285 277
2 1 27 0 0 4224 0 16 18 0 0 3
231 267
25 267
25 68
3 1 18 0 0 0 0 17 16 0 0 3
223 230
231 230
231 249
2 2 28 0 0 4224 0 18 17 0 0 3
19 68
19 239
174 239
3 1 19 0 0 0 0 21 17 0 0 4
171 194
176 194
176 221
174 221
3 2 29 0 0 4224 0 18 21 0 0 3
13 68
13 203
122 203
3 1 29 0 0 0 0 18 19 0 0 3
13 68
13 154
73 154
4 2 21 0 0 0 0 18 19 0 0 3
7 68
7 172
73 172
3 1 20 0 0 128 0 19 21 0 0 2
122 163
122 185
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
